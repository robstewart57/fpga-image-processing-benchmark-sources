-- ----------------------------------------------------------------------------
-- __  ___ __ ___  _ __   ___  ___ 
-- \ \/ / '__/ _ \| '_ \ / _ \/ __|
--  >  <| | | (_) | | | | (_) \__ \
-- /_/\_\_|  \___/|_| |_|\___/|___/
-- ----------------------------------------------------------------------------
-- Xronos synthesizer
-- Top level Network: ProgNetwork 
-- Date: 2017/11/02 14:01:53
-- ----------------------------------------------------------------------------

-- ----------------------------------------------------------------------------
-- Clock Domain(s) Information on the Network "ProgNetwork"
--
-- Network input port(s) clock domain:
--	In --> CLK
-- Network output port(s) clock domain:
-- 	Out --> CLK
-- 	dummy1 --> CLK
-- 	dummy2 --> CLK
-- 	dummy3 --> CLK
-- 	dummy4 --> CLK
-- Actor(s) clock domains:
--	LL1_H_iunzipFilter2D (LL1_H_iunzipFilter2D) --> CLK
--	HH1 (HH1) --> CLK
--	LL2_H_iunzipFilter2D (LL2_H_iunzipFilter2D) --> CLK
--	HH2 (HH2) --> CLK
--	LL3_H_iunzipFilter2D (LL3_H_iunzipFilter2D) --> CLK
--	HH3 (HH3) --> CLK
--	HL1 (HL1) --> CLK
--	HL2 (HL2) --> CLK
--	HL3 (HL3) --> CLK
--	LL1_L_iunzipFilter2D (LL1_L_iunzipFilter2D) --> CLK
--	LH1 (LH1) --> CLK
--	LL2_L_iunzipFilter2D (LL2_L_iunzipFilter2D) --> CLK
--	LH2 (LH2) --> CLK
--	LL3_L_iunzipFilter2D (LL3_L_iunzipFilter2D) --> CLK
--	LH3 (LH3) --> CLK
--	LL1 (LL1) --> CLK
--	image1_iunzip (image1_iunzip) --> CLK
--	LL1_H (LL1_H) --> CLK
--	LL1_L (LL1_L) --> CLK
--	LL2 (LL2) --> CLK
--	LL1_iunzip (LL1_iunzip) --> CLK
--	LL2_H (LL2_H) --> CLK
--	LL2_L (LL2_L) --> CLK
--	LL3 (LL3) --> CLK
--	LL2_iunzip (LL2_iunzip) --> CLK
--	LL3_H (LL3_H) --> CLK
--	LL3_L (LL3_L) --> CLK
--	image1 (image1) --> CLK
--	mapDia (mapDia) --> CLK
--	mapFinal (mapFinal) --> CLK
--	mapVer (mapVer) --> CLK
--	resized_HH1_xy (resized_HH1_xy) --> CLK
--	resized_HH1_xy_blurred (resized_HH1_xy_blurred) --> CLK
--	resized_HH2_xy (resized_HH2_xy) --> CLK
--	resized_HH2_xy_blurred (resized_HH2_xy_blurred) --> CLK
--	resized_HH3_xy (resized_HH3_xy) --> CLK
--	resized_HH3_xy_blurred (resized_HH3_xy_blurred) --> CLK
--	resized_LH1_xy (resized_LH1_xy) --> CLK
--	resized_LH1_xy_blurred (resized_LH1_xy_blurred) --> CLK
--	resized_LH2_xy (resized_LH2_xy) --> CLK
--	resized_LH2_xy_blurred (resized_LH2_xy_blurred) --> CLK
--	resized_LH3_xy (resized_LH3_xy) --> CLK
--	resized_LH3_xy_blurred (resized_LH3_xy_blurred) --> CLK

library ieee;
library SystemBuilder;

use ieee.std_logic_1164.all;

-- ----------------------------------------------------------------------------
-- Entity Declaration
-- ----------------------------------------------------------------------------
entity ProgNetwork is
port(
	 -- XDF Network Input(s)
	 In_data : in std_logic_vector(15 downto 0);
	 In_send : in std_logic;
	 In_ack : out std_logic;
	 In_rdy : out std_logic;
	 In_count : in std_logic_vector(15 downto 0);
	 -- XDF Network Output(s)
	 Out_data : out std_logic_vector(15 downto 0);
	 Out_send : out std_logic;
	 Out_ack : in std_logic;
	 Out_rdy : in std_logic;
	 Out_count : out std_logic_vector(15 downto 0);
	 dummy1_data : out std_logic_vector(15 downto 0);
	 dummy1_send : out std_logic;
	 dummy1_ack : in std_logic;
	 dummy1_rdy : in std_logic;
	 dummy1_count : out std_logic_vector(15 downto 0);
	 dummy2_data : out std_logic_vector(15 downto 0);
	 dummy2_send : out std_logic;
	 dummy2_ack : in std_logic;
	 dummy2_rdy : in std_logic;
	 dummy2_count : out std_logic_vector(15 downto 0);
	 dummy3_data : out std_logic_vector(15 downto 0);
	 dummy3_send : out std_logic;
	 dummy3_ack : in std_logic;
	 dummy3_rdy : in std_logic;
	 dummy3_count : out std_logic_vector(15 downto 0);
	 dummy4_data : out std_logic_vector(15 downto 0);
	 dummy4_send : out std_logic;
	 dummy4_ack : in std_logic;
	 dummy4_rdy : in std_logic;
	 dummy4_count : out std_logic_vector(15 downto 0);
	 -- Clock(s) and Reset
	 CLK : in std_logic;
	 RESET : in std_logic);
end entity ProgNetwork;

-- ----------------------------------------------------------------------------
-- Architecture Declaration
-- ----------------------------------------------------------------------------
architecture rtl of ProgNetwork is
	-- --------------------------------------------------------------------------
	-- Internal Signals
	-- --------------------------------------------------------------------------

	-- Clock(s) and Reset signal
	signal clocks, resets: std_logic_vector(0 downto 0);

	-- Network Input Port(s)
	signal ni_In_data : std_logic_vector(15 downto 0);
	signal ni_In_send : std_logic;
	signal ni_In_ack : std_logic;
	signal ni_In_rdy : std_logic;
	signal ni_In_count : std_logic_vector(15 downto 0);
	
	-- Network Input Port Fanout(s)
	signal nif_In_data : std_logic_vector(15 downto 0);
	signal nif_In_send : std_logic_vector(0 downto 0);
	signal nif_In_ack : std_logic_vector(0 downto 0);
	signal nif_In_rdy : std_logic_vector(0 downto 0);
	signal nif_In_count : std_logic_vector(15 downto 0);
	
	-- Network Output Port(s) 
	signal no_Out_data : std_logic_vector(15 downto 0);
	signal no_Out_send : std_logic;
	signal no_Out_ack : std_logic;
	signal no_Out_rdy : std_logic;
	signal no_Out_count : std_logic_vector(15 downto 0);
	signal no_dummy1_data : std_logic_vector(15 downto 0);
	signal no_dummy1_send : std_logic;
	signal no_dummy1_ack : std_logic;
	signal no_dummy1_rdy : std_logic;
	signal no_dummy1_count : std_logic_vector(15 downto 0);
	signal no_dummy2_data : std_logic_vector(15 downto 0);
	signal no_dummy2_send : std_logic;
	signal no_dummy2_ack : std_logic;
	signal no_dummy2_rdy : std_logic;
	signal no_dummy2_count : std_logic_vector(15 downto 0);
	signal no_dummy3_data : std_logic_vector(15 downto 0);
	signal no_dummy3_send : std_logic;
	signal no_dummy3_ack : std_logic;
	signal no_dummy3_rdy : std_logic;
	signal no_dummy3_count : std_logic_vector(15 downto 0);
	signal no_dummy4_data : std_logic_vector(15 downto 0);
	signal no_dummy4_send : std_logic;
	signal no_dummy4_ack : std_logic;
	signal no_dummy4_rdy : std_logic;
	signal no_dummy4_count : std_logic_vector(15 downto 0);
	
	-- Actors Input/Output and Output fanout signals
	signal ai_LL1_H_iunzipFilter2D_In1_data : std_logic_vector(15 downto 0);
	signal ai_LL1_H_iunzipFilter2D_In1_send : std_logic;
	signal ai_LL1_H_iunzipFilter2D_In1_ack : std_logic;
	signal ai_LL1_H_iunzipFilter2D_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_LL1_H_iunzipFilter2D_Out1_data : std_logic_vector(15 downto 0);
	signal ao_LL1_H_iunzipFilter2D_Out1_send : std_logic;
	signal ao_LL1_H_iunzipFilter2D_Out1_ack : std_logic;
	signal ao_LL1_H_iunzipFilter2D_Out1_rdy : std_logic;
	signal ao_LL1_H_iunzipFilter2D_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_LL1_H_iunzipFilter2D_Out1_data : std_logic_vector(15 downto 0);
	signal aof_LL1_H_iunzipFilter2D_Out1_send : std_logic_vector(0 downto 0);
	signal aof_LL1_H_iunzipFilter2D_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_LL1_H_iunzipFilter2D_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_LL1_H_iunzipFilter2D_Out1_count : std_logic_vector(15 downto 0);
	
	signal ao_LL1_H_iunzipFilter2D_Out2_data : std_logic_vector(15 downto 0);
	signal ao_LL1_H_iunzipFilter2D_Out2_send : std_logic;
	signal ao_LL1_H_iunzipFilter2D_Out2_ack : std_logic;
	signal ao_LL1_H_iunzipFilter2D_Out2_rdy : std_logic;
	signal ao_LL1_H_iunzipFilter2D_Out2_count : std_logic_vector(15 downto 0);
	
	signal aof_LL1_H_iunzipFilter2D_Out2_data : std_logic_vector(15 downto 0);
	signal aof_LL1_H_iunzipFilter2D_Out2_send : std_logic_vector(0 downto 0);
	signal aof_LL1_H_iunzipFilter2D_Out2_ack : std_logic_vector(0 downto 0);
	signal aof_LL1_H_iunzipFilter2D_Out2_rdy : std_logic_vector(0 downto 0);
	signal aof_LL1_H_iunzipFilter2D_Out2_count : std_logic_vector(15 downto 0);
	
	signal ai_HH1_In1_data : std_logic_vector(15 downto 0);
	signal ai_HH1_In1_send : std_logic;
	signal ai_HH1_In1_ack : std_logic;
	signal ai_HH1_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_HH1_Out1_data : std_logic_vector(15 downto 0);
	signal ao_HH1_Out1_send : std_logic;
	signal ao_HH1_Out1_ack : std_logic;
	signal ao_HH1_Out1_rdy : std_logic;
	signal ao_HH1_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_HH1_Out1_data : std_logic_vector(15 downto 0);
	signal aof_HH1_Out1_send : std_logic_vector(0 downto 0);
	signal aof_HH1_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_HH1_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_HH1_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_LL2_H_iunzipFilter2D_In1_data : std_logic_vector(15 downto 0);
	signal ai_LL2_H_iunzipFilter2D_In1_send : std_logic;
	signal ai_LL2_H_iunzipFilter2D_In1_ack : std_logic;
	signal ai_LL2_H_iunzipFilter2D_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_LL2_H_iunzipFilter2D_Out1_data : std_logic_vector(15 downto 0);
	signal ao_LL2_H_iunzipFilter2D_Out1_send : std_logic;
	signal ao_LL2_H_iunzipFilter2D_Out1_ack : std_logic;
	signal ao_LL2_H_iunzipFilter2D_Out1_rdy : std_logic;
	signal ao_LL2_H_iunzipFilter2D_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_LL2_H_iunzipFilter2D_Out1_data : std_logic_vector(15 downto 0);
	signal aof_LL2_H_iunzipFilter2D_Out1_send : std_logic_vector(0 downto 0);
	signal aof_LL2_H_iunzipFilter2D_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_LL2_H_iunzipFilter2D_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_LL2_H_iunzipFilter2D_Out1_count : std_logic_vector(15 downto 0);
	
	signal ao_LL2_H_iunzipFilter2D_Out2_data : std_logic_vector(15 downto 0);
	signal ao_LL2_H_iunzipFilter2D_Out2_send : std_logic;
	signal ao_LL2_H_iunzipFilter2D_Out2_ack : std_logic;
	signal ao_LL2_H_iunzipFilter2D_Out2_rdy : std_logic;
	signal ao_LL2_H_iunzipFilter2D_Out2_count : std_logic_vector(15 downto 0);
	
	signal aof_LL2_H_iunzipFilter2D_Out2_data : std_logic_vector(15 downto 0);
	signal aof_LL2_H_iunzipFilter2D_Out2_send : std_logic_vector(0 downto 0);
	signal aof_LL2_H_iunzipFilter2D_Out2_ack : std_logic_vector(0 downto 0);
	signal aof_LL2_H_iunzipFilter2D_Out2_rdy : std_logic_vector(0 downto 0);
	signal aof_LL2_H_iunzipFilter2D_Out2_count : std_logic_vector(15 downto 0);
	
	signal ai_HH2_In1_data : std_logic_vector(15 downto 0);
	signal ai_HH2_In1_send : std_logic;
	signal ai_HH2_In1_ack : std_logic;
	signal ai_HH2_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_HH2_Out1_data : std_logic_vector(15 downto 0);
	signal ao_HH2_Out1_send : std_logic;
	signal ao_HH2_Out1_ack : std_logic;
	signal ao_HH2_Out1_rdy : std_logic;
	signal ao_HH2_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_HH2_Out1_data : std_logic_vector(15 downto 0);
	signal aof_HH2_Out1_send : std_logic_vector(0 downto 0);
	signal aof_HH2_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_HH2_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_HH2_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_LL3_H_iunzipFilter2D_In1_data : std_logic_vector(15 downto 0);
	signal ai_LL3_H_iunzipFilter2D_In1_send : std_logic;
	signal ai_LL3_H_iunzipFilter2D_In1_ack : std_logic;
	signal ai_LL3_H_iunzipFilter2D_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_LL3_H_iunzipFilter2D_Out1_data : std_logic_vector(15 downto 0);
	signal ao_LL3_H_iunzipFilter2D_Out1_send : std_logic;
	signal ao_LL3_H_iunzipFilter2D_Out1_ack : std_logic;
	signal ao_LL3_H_iunzipFilter2D_Out1_rdy : std_logic;
	signal ao_LL3_H_iunzipFilter2D_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_LL3_H_iunzipFilter2D_Out1_data : std_logic_vector(15 downto 0);
	signal aof_LL3_H_iunzipFilter2D_Out1_send : std_logic_vector(0 downto 0);
	signal aof_LL3_H_iunzipFilter2D_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_LL3_H_iunzipFilter2D_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_LL3_H_iunzipFilter2D_Out1_count : std_logic_vector(15 downto 0);
	
	signal ao_LL3_H_iunzipFilter2D_Out2_data : std_logic_vector(15 downto 0);
	signal ao_LL3_H_iunzipFilter2D_Out2_send : std_logic;
	signal ao_LL3_H_iunzipFilter2D_Out2_ack : std_logic;
	signal ao_LL3_H_iunzipFilter2D_Out2_rdy : std_logic;
	signal ao_LL3_H_iunzipFilter2D_Out2_count : std_logic_vector(15 downto 0);
	
	signal aof_LL3_H_iunzipFilter2D_Out2_data : std_logic_vector(15 downto 0);
	signal aof_LL3_H_iunzipFilter2D_Out2_send : std_logic_vector(0 downto 0);
	signal aof_LL3_H_iunzipFilter2D_Out2_ack : std_logic_vector(0 downto 0);
	signal aof_LL3_H_iunzipFilter2D_Out2_rdy : std_logic_vector(0 downto 0);
	signal aof_LL3_H_iunzipFilter2D_Out2_count : std_logic_vector(15 downto 0);
	
	signal ai_HH3_In1_data : std_logic_vector(15 downto 0);
	signal ai_HH3_In1_send : std_logic;
	signal ai_HH3_In1_ack : std_logic;
	signal ai_HH3_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_HH3_Out1_data : std_logic_vector(15 downto 0);
	signal ao_HH3_Out1_send : std_logic;
	signal ao_HH3_Out1_ack : std_logic;
	signal ao_HH3_Out1_rdy : std_logic;
	signal ao_HH3_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_HH3_Out1_data : std_logic_vector(15 downto 0);
	signal aof_HH3_Out1_send : std_logic_vector(0 downto 0);
	signal aof_HH3_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_HH3_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_HH3_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_HL1_In1_data : std_logic_vector(15 downto 0);
	signal ai_HL1_In1_send : std_logic;
	signal ai_HL1_In1_ack : std_logic;
	signal ai_HL1_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_HL1_Out1_data : std_logic_vector(15 downto 0);
	signal ao_HL1_Out1_send : std_logic;
	signal ao_HL1_Out1_ack : std_logic;
	signal ao_HL1_Out1_rdy : std_logic;
	signal ao_HL1_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_HL1_Out1_data : std_logic_vector(15 downto 0);
	signal aof_HL1_Out1_send : std_logic_vector(0 downto 0);
	signal aof_HL1_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_HL1_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_HL1_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_HL2_In1_data : std_logic_vector(15 downto 0);
	signal ai_HL2_In1_send : std_logic;
	signal ai_HL2_In1_ack : std_logic;
	signal ai_HL2_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_HL2_Out1_data : std_logic_vector(15 downto 0);
	signal ao_HL2_Out1_send : std_logic;
	signal ao_HL2_Out1_ack : std_logic;
	signal ao_HL2_Out1_rdy : std_logic;
	signal ao_HL2_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_HL2_Out1_data : std_logic_vector(15 downto 0);
	signal aof_HL2_Out1_send : std_logic_vector(0 downto 0);
	signal aof_HL2_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_HL2_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_HL2_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_HL3_In1_data : std_logic_vector(15 downto 0);
	signal ai_HL3_In1_send : std_logic;
	signal ai_HL3_In1_ack : std_logic;
	signal ai_HL3_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_HL3_Out1_data : std_logic_vector(15 downto 0);
	signal ao_HL3_Out1_send : std_logic;
	signal ao_HL3_Out1_ack : std_logic;
	signal ao_HL3_Out1_rdy : std_logic;
	signal ao_HL3_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_HL3_Out1_data : std_logic_vector(15 downto 0);
	signal aof_HL3_Out1_send : std_logic_vector(0 downto 0);
	signal aof_HL3_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_HL3_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_HL3_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_LL1_L_iunzipFilter2D_In1_data : std_logic_vector(15 downto 0);
	signal ai_LL1_L_iunzipFilter2D_In1_send : std_logic;
	signal ai_LL1_L_iunzipFilter2D_In1_ack : std_logic;
	signal ai_LL1_L_iunzipFilter2D_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_LL1_L_iunzipFilter2D_Out1_data : std_logic_vector(15 downto 0);
	signal ao_LL1_L_iunzipFilter2D_Out1_send : std_logic;
	signal ao_LL1_L_iunzipFilter2D_Out1_ack : std_logic;
	signal ao_LL1_L_iunzipFilter2D_Out1_rdy : std_logic;
	signal ao_LL1_L_iunzipFilter2D_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_LL1_L_iunzipFilter2D_Out1_data : std_logic_vector(15 downto 0);
	signal aof_LL1_L_iunzipFilter2D_Out1_send : std_logic_vector(0 downto 0);
	signal aof_LL1_L_iunzipFilter2D_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_LL1_L_iunzipFilter2D_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_LL1_L_iunzipFilter2D_Out1_count : std_logic_vector(15 downto 0);
	
	signal ao_LL1_L_iunzipFilter2D_Out2_data : std_logic_vector(15 downto 0);
	signal ao_LL1_L_iunzipFilter2D_Out2_send : std_logic;
	signal ao_LL1_L_iunzipFilter2D_Out2_ack : std_logic;
	signal ao_LL1_L_iunzipFilter2D_Out2_rdy : std_logic;
	signal ao_LL1_L_iunzipFilter2D_Out2_count : std_logic_vector(15 downto 0);
	
	signal aof_LL1_L_iunzipFilter2D_Out2_data : std_logic_vector(15 downto 0);
	signal aof_LL1_L_iunzipFilter2D_Out2_send : std_logic_vector(0 downto 0);
	signal aof_LL1_L_iunzipFilter2D_Out2_ack : std_logic_vector(0 downto 0);
	signal aof_LL1_L_iunzipFilter2D_Out2_rdy : std_logic_vector(0 downto 0);
	signal aof_LL1_L_iunzipFilter2D_Out2_count : std_logic_vector(15 downto 0);
	
	signal ai_LH1_In1_data : std_logic_vector(15 downto 0);
	signal ai_LH1_In1_send : std_logic;
	signal ai_LH1_In1_ack : std_logic;
	signal ai_LH1_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_LH1_Out1_data : std_logic_vector(15 downto 0);
	signal ao_LH1_Out1_send : std_logic;
	signal ao_LH1_Out1_ack : std_logic;
	signal ao_LH1_Out1_rdy : std_logic;
	signal ao_LH1_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_LH1_Out1_data : std_logic_vector(15 downto 0);
	signal aof_LH1_Out1_send : std_logic_vector(0 downto 0);
	signal aof_LH1_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_LH1_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_LH1_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_LL2_L_iunzipFilter2D_In1_data : std_logic_vector(15 downto 0);
	signal ai_LL2_L_iunzipFilter2D_In1_send : std_logic;
	signal ai_LL2_L_iunzipFilter2D_In1_ack : std_logic;
	signal ai_LL2_L_iunzipFilter2D_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_LL2_L_iunzipFilter2D_Out1_data : std_logic_vector(15 downto 0);
	signal ao_LL2_L_iunzipFilter2D_Out1_send : std_logic;
	signal ao_LL2_L_iunzipFilter2D_Out1_ack : std_logic;
	signal ao_LL2_L_iunzipFilter2D_Out1_rdy : std_logic;
	signal ao_LL2_L_iunzipFilter2D_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_LL2_L_iunzipFilter2D_Out1_data : std_logic_vector(15 downto 0);
	signal aof_LL2_L_iunzipFilter2D_Out1_send : std_logic_vector(0 downto 0);
	signal aof_LL2_L_iunzipFilter2D_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_LL2_L_iunzipFilter2D_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_LL2_L_iunzipFilter2D_Out1_count : std_logic_vector(15 downto 0);
	
	signal ao_LL2_L_iunzipFilter2D_Out2_data : std_logic_vector(15 downto 0);
	signal ao_LL2_L_iunzipFilter2D_Out2_send : std_logic;
	signal ao_LL2_L_iunzipFilter2D_Out2_ack : std_logic;
	signal ao_LL2_L_iunzipFilter2D_Out2_rdy : std_logic;
	signal ao_LL2_L_iunzipFilter2D_Out2_count : std_logic_vector(15 downto 0);
	
	signal aof_LL2_L_iunzipFilter2D_Out2_data : std_logic_vector(15 downto 0);
	signal aof_LL2_L_iunzipFilter2D_Out2_send : std_logic_vector(0 downto 0);
	signal aof_LL2_L_iunzipFilter2D_Out2_ack : std_logic_vector(0 downto 0);
	signal aof_LL2_L_iunzipFilter2D_Out2_rdy : std_logic_vector(0 downto 0);
	signal aof_LL2_L_iunzipFilter2D_Out2_count : std_logic_vector(15 downto 0);
	
	signal ai_LH2_In1_data : std_logic_vector(15 downto 0);
	signal ai_LH2_In1_send : std_logic;
	signal ai_LH2_In1_ack : std_logic;
	signal ai_LH2_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_LH2_Out1_data : std_logic_vector(15 downto 0);
	signal ao_LH2_Out1_send : std_logic;
	signal ao_LH2_Out1_ack : std_logic;
	signal ao_LH2_Out1_rdy : std_logic;
	signal ao_LH2_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_LH2_Out1_data : std_logic_vector(15 downto 0);
	signal aof_LH2_Out1_send : std_logic_vector(0 downto 0);
	signal aof_LH2_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_LH2_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_LH2_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_LL3_L_iunzipFilter2D_In1_data : std_logic_vector(15 downto 0);
	signal ai_LL3_L_iunzipFilter2D_In1_send : std_logic;
	signal ai_LL3_L_iunzipFilter2D_In1_ack : std_logic;
	signal ai_LL3_L_iunzipFilter2D_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_LL3_L_iunzipFilter2D_Out1_data : std_logic_vector(15 downto 0);
	signal ao_LL3_L_iunzipFilter2D_Out1_send : std_logic;
	signal ao_LL3_L_iunzipFilter2D_Out1_ack : std_logic;
	signal ao_LL3_L_iunzipFilter2D_Out1_rdy : std_logic;
	signal ao_LL3_L_iunzipFilter2D_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_LL3_L_iunzipFilter2D_Out1_data : std_logic_vector(15 downto 0);
	signal aof_LL3_L_iunzipFilter2D_Out1_send : std_logic_vector(0 downto 0);
	signal aof_LL3_L_iunzipFilter2D_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_LL3_L_iunzipFilter2D_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_LL3_L_iunzipFilter2D_Out1_count : std_logic_vector(15 downto 0);
	
	signal ao_LL3_L_iunzipFilter2D_Out2_data : std_logic_vector(15 downto 0);
	signal ao_LL3_L_iunzipFilter2D_Out2_send : std_logic;
	signal ao_LL3_L_iunzipFilter2D_Out2_ack : std_logic;
	signal ao_LL3_L_iunzipFilter2D_Out2_rdy : std_logic;
	signal ao_LL3_L_iunzipFilter2D_Out2_count : std_logic_vector(15 downto 0);
	
	signal aof_LL3_L_iunzipFilter2D_Out2_data : std_logic_vector(15 downto 0);
	signal aof_LL3_L_iunzipFilter2D_Out2_send : std_logic_vector(0 downto 0);
	signal aof_LL3_L_iunzipFilter2D_Out2_ack : std_logic_vector(0 downto 0);
	signal aof_LL3_L_iunzipFilter2D_Out2_rdy : std_logic_vector(0 downto 0);
	signal aof_LL3_L_iunzipFilter2D_Out2_count : std_logic_vector(15 downto 0);
	
	signal ai_LH3_In1_data : std_logic_vector(15 downto 0);
	signal ai_LH3_In1_send : std_logic;
	signal ai_LH3_In1_ack : std_logic;
	signal ai_LH3_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_LH3_Out1_data : std_logic_vector(15 downto 0);
	signal ao_LH3_Out1_send : std_logic;
	signal ao_LH3_Out1_ack : std_logic;
	signal ao_LH3_Out1_rdy : std_logic;
	signal ao_LH3_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_LH3_Out1_data : std_logic_vector(15 downto 0);
	signal aof_LH3_Out1_send : std_logic_vector(0 downto 0);
	signal aof_LH3_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_LH3_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_LH3_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_LL1_In1_data : std_logic_vector(15 downto 0);
	signal ai_LL1_In1_send : std_logic;
	signal ai_LL1_In1_ack : std_logic;
	signal ai_LL1_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_LL1_Out1_data : std_logic_vector(15 downto 0);
	signal ao_LL1_Out1_send : std_logic;
	signal ao_LL1_Out1_ack : std_logic;
	signal ao_LL1_Out1_rdy : std_logic;
	signal ao_LL1_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_LL1_Out1_data : std_logic_vector(15 downto 0);
	signal aof_LL1_Out1_send : std_logic_vector(0 downto 0);
	signal aof_LL1_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_LL1_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_LL1_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_image1_iunzip_In1_data : std_logic_vector(15 downto 0);
	signal ai_image1_iunzip_In1_send : std_logic;
	signal ai_image1_iunzip_In1_ack : std_logic;
	signal ai_image1_iunzip_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_image1_iunzip_Out1_data : std_logic_vector(15 downto 0);
	signal ao_image1_iunzip_Out1_send : std_logic;
	signal ao_image1_iunzip_Out1_ack : std_logic;
	signal ao_image1_iunzip_Out1_rdy : std_logic;
	signal ao_image1_iunzip_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_image1_iunzip_Out1_data : std_logic_vector(15 downto 0);
	signal aof_image1_iunzip_Out1_send : std_logic_vector(0 downto 0);
	signal aof_image1_iunzip_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_image1_iunzip_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_image1_iunzip_Out1_count : std_logic_vector(15 downto 0);
	
	signal ao_image1_iunzip_Out2_data : std_logic_vector(15 downto 0);
	signal ao_image1_iunzip_Out2_send : std_logic;
	signal ao_image1_iunzip_Out2_ack : std_logic;
	signal ao_image1_iunzip_Out2_rdy : std_logic;
	signal ao_image1_iunzip_Out2_count : std_logic_vector(15 downto 0);
	
	signal aof_image1_iunzip_Out2_data : std_logic_vector(15 downto 0);
	signal aof_image1_iunzip_Out2_send : std_logic_vector(0 downto 0);
	signal aof_image1_iunzip_Out2_ack : std_logic_vector(0 downto 0);
	signal aof_image1_iunzip_Out2_rdy : std_logic_vector(0 downto 0);
	signal aof_image1_iunzip_Out2_count : std_logic_vector(15 downto 0);
	
	signal ai_LL1_H_In1_data : std_logic_vector(15 downto 0);
	signal ai_LL1_H_In1_send : std_logic;
	signal ai_LL1_H_In1_ack : std_logic;
	signal ai_LL1_H_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_LL1_H_Out1_data : std_logic_vector(15 downto 0);
	signal ao_LL1_H_Out1_send : std_logic;
	signal ao_LL1_H_Out1_ack : std_logic;
	signal ao_LL1_H_Out1_rdy : std_logic;
	signal ao_LL1_H_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_LL1_H_Out1_data : std_logic_vector(15 downto 0);
	signal aof_LL1_H_Out1_send : std_logic_vector(0 downto 0);
	signal aof_LL1_H_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_LL1_H_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_LL1_H_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_LL1_L_In1_data : std_logic_vector(15 downto 0);
	signal ai_LL1_L_In1_send : std_logic;
	signal ai_LL1_L_In1_ack : std_logic;
	signal ai_LL1_L_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_LL1_L_Out1_data : std_logic_vector(15 downto 0);
	signal ao_LL1_L_Out1_send : std_logic;
	signal ao_LL1_L_Out1_ack : std_logic;
	signal ao_LL1_L_Out1_rdy : std_logic;
	signal ao_LL1_L_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_LL1_L_Out1_data : std_logic_vector(15 downto 0);
	signal aof_LL1_L_Out1_send : std_logic_vector(0 downto 0);
	signal aof_LL1_L_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_LL1_L_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_LL1_L_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_LL2_In1_data : std_logic_vector(15 downto 0);
	signal ai_LL2_In1_send : std_logic;
	signal ai_LL2_In1_ack : std_logic;
	signal ai_LL2_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_LL2_Out1_data : std_logic_vector(15 downto 0);
	signal ao_LL2_Out1_send : std_logic;
	signal ao_LL2_Out1_ack : std_logic;
	signal ao_LL2_Out1_rdy : std_logic;
	signal ao_LL2_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_LL2_Out1_data : std_logic_vector(15 downto 0);
	signal aof_LL2_Out1_send : std_logic_vector(0 downto 0);
	signal aof_LL2_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_LL2_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_LL2_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_LL1_iunzip_In1_data : std_logic_vector(15 downto 0);
	signal ai_LL1_iunzip_In1_send : std_logic;
	signal ai_LL1_iunzip_In1_ack : std_logic;
	signal ai_LL1_iunzip_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_LL1_iunzip_Out1_data : std_logic_vector(15 downto 0);
	signal ao_LL1_iunzip_Out1_send : std_logic;
	signal ao_LL1_iunzip_Out1_ack : std_logic;
	signal ao_LL1_iunzip_Out1_rdy : std_logic;
	signal ao_LL1_iunzip_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_LL1_iunzip_Out1_data : std_logic_vector(15 downto 0);
	signal aof_LL1_iunzip_Out1_send : std_logic_vector(0 downto 0);
	signal aof_LL1_iunzip_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_LL1_iunzip_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_LL1_iunzip_Out1_count : std_logic_vector(15 downto 0);
	
	signal ao_LL1_iunzip_Out2_data : std_logic_vector(15 downto 0);
	signal ao_LL1_iunzip_Out2_send : std_logic;
	signal ao_LL1_iunzip_Out2_ack : std_logic;
	signal ao_LL1_iunzip_Out2_rdy : std_logic;
	signal ao_LL1_iunzip_Out2_count : std_logic_vector(15 downto 0);
	
	signal aof_LL1_iunzip_Out2_data : std_logic_vector(15 downto 0);
	signal aof_LL1_iunzip_Out2_send : std_logic_vector(0 downto 0);
	signal aof_LL1_iunzip_Out2_ack : std_logic_vector(0 downto 0);
	signal aof_LL1_iunzip_Out2_rdy : std_logic_vector(0 downto 0);
	signal aof_LL1_iunzip_Out2_count : std_logic_vector(15 downto 0);
	
	signal ai_LL2_H_In1_data : std_logic_vector(15 downto 0);
	signal ai_LL2_H_In1_send : std_logic;
	signal ai_LL2_H_In1_ack : std_logic;
	signal ai_LL2_H_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_LL2_H_Out1_data : std_logic_vector(15 downto 0);
	signal ao_LL2_H_Out1_send : std_logic;
	signal ao_LL2_H_Out1_ack : std_logic;
	signal ao_LL2_H_Out1_rdy : std_logic;
	signal ao_LL2_H_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_LL2_H_Out1_data : std_logic_vector(15 downto 0);
	signal aof_LL2_H_Out1_send : std_logic_vector(0 downto 0);
	signal aof_LL2_H_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_LL2_H_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_LL2_H_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_LL2_L_In1_data : std_logic_vector(15 downto 0);
	signal ai_LL2_L_In1_send : std_logic;
	signal ai_LL2_L_In1_ack : std_logic;
	signal ai_LL2_L_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_LL2_L_Out1_data : std_logic_vector(15 downto 0);
	signal ao_LL2_L_Out1_send : std_logic;
	signal ao_LL2_L_Out1_ack : std_logic;
	signal ao_LL2_L_Out1_rdy : std_logic;
	signal ao_LL2_L_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_LL2_L_Out1_data : std_logic_vector(15 downto 0);
	signal aof_LL2_L_Out1_send : std_logic_vector(0 downto 0);
	signal aof_LL2_L_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_LL2_L_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_LL2_L_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_LL3_In1_data : std_logic_vector(15 downto 0);
	signal ai_LL3_In1_send : std_logic;
	signal ai_LL3_In1_ack : std_logic;
	signal ai_LL3_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_LL3_Out1_data : std_logic_vector(15 downto 0);
	signal ao_LL3_Out1_send : std_logic;
	signal ao_LL3_Out1_ack : std_logic;
	signal ao_LL3_Out1_rdy : std_logic;
	signal ao_LL3_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_LL3_Out1_data : std_logic_vector(15 downto 0);
	signal aof_LL3_Out1_send : std_logic_vector(0 downto 0);
	signal aof_LL3_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_LL3_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_LL3_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_LL2_iunzip_In1_data : std_logic_vector(15 downto 0);
	signal ai_LL2_iunzip_In1_send : std_logic;
	signal ai_LL2_iunzip_In1_ack : std_logic;
	signal ai_LL2_iunzip_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_LL2_iunzip_Out1_data : std_logic_vector(15 downto 0);
	signal ao_LL2_iunzip_Out1_send : std_logic;
	signal ao_LL2_iunzip_Out1_ack : std_logic;
	signal ao_LL2_iunzip_Out1_rdy : std_logic;
	signal ao_LL2_iunzip_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_LL2_iunzip_Out1_data : std_logic_vector(15 downto 0);
	signal aof_LL2_iunzip_Out1_send : std_logic_vector(0 downto 0);
	signal aof_LL2_iunzip_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_LL2_iunzip_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_LL2_iunzip_Out1_count : std_logic_vector(15 downto 0);
	
	signal ao_LL2_iunzip_Out2_data : std_logic_vector(15 downto 0);
	signal ao_LL2_iunzip_Out2_send : std_logic;
	signal ao_LL2_iunzip_Out2_ack : std_logic;
	signal ao_LL2_iunzip_Out2_rdy : std_logic;
	signal ao_LL2_iunzip_Out2_count : std_logic_vector(15 downto 0);
	
	signal aof_LL2_iunzip_Out2_data : std_logic_vector(15 downto 0);
	signal aof_LL2_iunzip_Out2_send : std_logic_vector(0 downto 0);
	signal aof_LL2_iunzip_Out2_ack : std_logic_vector(0 downto 0);
	signal aof_LL2_iunzip_Out2_rdy : std_logic_vector(0 downto 0);
	signal aof_LL2_iunzip_Out2_count : std_logic_vector(15 downto 0);
	
	signal ai_LL3_H_In1_data : std_logic_vector(15 downto 0);
	signal ai_LL3_H_In1_send : std_logic;
	signal ai_LL3_H_In1_ack : std_logic;
	signal ai_LL3_H_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_LL3_H_Out1_data : std_logic_vector(15 downto 0);
	signal ao_LL3_H_Out1_send : std_logic;
	signal ao_LL3_H_Out1_ack : std_logic;
	signal ao_LL3_H_Out1_rdy : std_logic;
	signal ao_LL3_H_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_LL3_H_Out1_data : std_logic_vector(15 downto 0);
	signal aof_LL3_H_Out1_send : std_logic_vector(0 downto 0);
	signal aof_LL3_H_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_LL3_H_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_LL3_H_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_LL3_L_In1_data : std_logic_vector(15 downto 0);
	signal ai_LL3_L_In1_send : std_logic;
	signal ai_LL3_L_In1_ack : std_logic;
	signal ai_LL3_L_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_LL3_L_Out1_data : std_logic_vector(15 downto 0);
	signal ao_LL3_L_Out1_send : std_logic;
	signal ao_LL3_L_Out1_ack : std_logic;
	signal ao_LL3_L_Out1_rdy : std_logic;
	signal ao_LL3_L_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_LL3_L_Out1_data : std_logic_vector(15 downto 0);
	signal aof_LL3_L_Out1_send : std_logic_vector(0 downto 0);
	signal aof_LL3_L_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_LL3_L_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_LL3_L_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_image1_In1_data : std_logic_vector(15 downto 0);
	signal ai_image1_In1_send : std_logic;
	signal ai_image1_In1_ack : std_logic;
	signal ai_image1_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_image1_Out1_data : std_logic_vector(15 downto 0);
	signal ao_image1_Out1_send : std_logic;
	signal ao_image1_Out1_ack : std_logic;
	signal ao_image1_Out1_rdy : std_logic;
	signal ao_image1_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_image1_Out1_data : std_logic_vector(15 downto 0);
	signal aof_image1_Out1_send : std_logic_vector(0 downto 0);
	signal aof_image1_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_image1_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_image1_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_mapDia_In1_data : std_logic_vector(15 downto 0);
	signal ai_mapDia_In1_send : std_logic;
	signal ai_mapDia_In1_ack : std_logic;
	signal ai_mapDia_In1_count : std_logic_vector(15 downto 0);
	
	signal ai_mapDia_In2_data : std_logic_vector(15 downto 0);
	signal ai_mapDia_In2_send : std_logic;
	signal ai_mapDia_In2_ack : std_logic;
	signal ai_mapDia_In2_count : std_logic_vector(15 downto 0);
	
	signal ai_mapDia_In3_data : std_logic_vector(15 downto 0);
	signal ai_mapDia_In3_send : std_logic;
	signal ai_mapDia_In3_ack : std_logic;
	signal ai_mapDia_In3_count : std_logic_vector(15 downto 0);
	
	signal ao_mapDia_Out1_data : std_logic_vector(15 downto 0);
	signal ao_mapDia_Out1_send : std_logic;
	signal ao_mapDia_Out1_ack : std_logic;
	signal ao_mapDia_Out1_rdy : std_logic;
	signal ao_mapDia_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_mapDia_Out1_data : std_logic_vector(15 downto 0);
	signal aof_mapDia_Out1_send : std_logic_vector(0 downto 0);
	signal aof_mapDia_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_mapDia_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_mapDia_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_mapFinal_In1_data : std_logic_vector(15 downto 0);
	signal ai_mapFinal_In1_send : std_logic;
	signal ai_mapFinal_In1_ack : std_logic;
	signal ai_mapFinal_In1_count : std_logic_vector(15 downto 0);
	
	signal ai_mapFinal_In2_data : std_logic_vector(15 downto 0);
	signal ai_mapFinal_In2_send : std_logic;
	signal ai_mapFinal_In2_ack : std_logic;
	signal ai_mapFinal_In2_count : std_logic_vector(15 downto 0);
	
	signal ao_mapFinal_Out1_data : std_logic_vector(15 downto 0);
	signal ao_mapFinal_Out1_send : std_logic;
	signal ao_mapFinal_Out1_ack : std_logic;
	signal ao_mapFinal_Out1_rdy : std_logic;
	signal ao_mapFinal_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_mapFinal_Out1_data : std_logic_vector(15 downto 0);
	signal aof_mapFinal_Out1_send : std_logic_vector(0 downto 0);
	signal aof_mapFinal_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_mapFinal_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_mapFinal_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_mapVer_In1_data : std_logic_vector(15 downto 0);
	signal ai_mapVer_In1_send : std_logic;
	signal ai_mapVer_In1_ack : std_logic;
	signal ai_mapVer_In1_count : std_logic_vector(15 downto 0);
	
	signal ai_mapVer_In2_data : std_logic_vector(15 downto 0);
	signal ai_mapVer_In2_send : std_logic;
	signal ai_mapVer_In2_ack : std_logic;
	signal ai_mapVer_In2_count : std_logic_vector(15 downto 0);
	
	signal ai_mapVer_In3_data : std_logic_vector(15 downto 0);
	signal ai_mapVer_In3_send : std_logic;
	signal ai_mapVer_In3_ack : std_logic;
	signal ai_mapVer_In3_count : std_logic_vector(15 downto 0);
	
	signal ao_mapVer_Out1_data : std_logic_vector(15 downto 0);
	signal ao_mapVer_Out1_send : std_logic;
	signal ao_mapVer_Out1_ack : std_logic;
	signal ao_mapVer_Out1_rdy : std_logic;
	signal ao_mapVer_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_mapVer_Out1_data : std_logic_vector(15 downto 0);
	signal aof_mapVer_Out1_send : std_logic_vector(0 downto 0);
	signal aof_mapVer_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_mapVer_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_mapVer_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_resized_HH1_xy_In1_data : std_logic_vector(15 downto 0);
	signal ai_resized_HH1_xy_In1_send : std_logic;
	signal ai_resized_HH1_xy_In1_ack : std_logic;
	signal ai_resized_HH1_xy_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_resized_HH1_xy_Out1_data : std_logic_vector(15 downto 0);
	signal ao_resized_HH1_xy_Out1_send : std_logic;
	signal ao_resized_HH1_xy_Out1_ack : std_logic;
	signal ao_resized_HH1_xy_Out1_rdy : std_logic;
	signal ao_resized_HH1_xy_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_resized_HH1_xy_Out1_data : std_logic_vector(15 downto 0);
	signal aof_resized_HH1_xy_Out1_send : std_logic_vector(0 downto 0);
	signal aof_resized_HH1_xy_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_resized_HH1_xy_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_resized_HH1_xy_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_resized_HH1_xy_blurred_In1_data : std_logic_vector(15 downto 0);
	signal ai_resized_HH1_xy_blurred_In1_send : std_logic;
	signal ai_resized_HH1_xy_blurred_In1_ack : std_logic;
	signal ai_resized_HH1_xy_blurred_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_resized_HH1_xy_blurred_Out1_data : std_logic_vector(15 downto 0);
	signal ao_resized_HH1_xy_blurred_Out1_send : std_logic;
	signal ao_resized_HH1_xy_blurred_Out1_ack : std_logic;
	signal ao_resized_HH1_xy_blurred_Out1_rdy : std_logic;
	signal ao_resized_HH1_xy_blurred_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_resized_HH1_xy_blurred_Out1_data : std_logic_vector(15 downto 0);
	signal aof_resized_HH1_xy_blurred_Out1_send : std_logic_vector(0 downto 0);
	signal aof_resized_HH1_xy_blurred_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_resized_HH1_xy_blurred_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_resized_HH1_xy_blurred_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_resized_HH2_xy_In1_data : std_logic_vector(15 downto 0);
	signal ai_resized_HH2_xy_In1_send : std_logic;
	signal ai_resized_HH2_xy_In1_ack : std_logic;
	signal ai_resized_HH2_xy_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_resized_HH2_xy_Out1_data : std_logic_vector(15 downto 0);
	signal ao_resized_HH2_xy_Out1_send : std_logic;
	signal ao_resized_HH2_xy_Out1_ack : std_logic;
	signal ao_resized_HH2_xy_Out1_rdy : std_logic;
	signal ao_resized_HH2_xy_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_resized_HH2_xy_Out1_data : std_logic_vector(15 downto 0);
	signal aof_resized_HH2_xy_Out1_send : std_logic_vector(0 downto 0);
	signal aof_resized_HH2_xy_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_resized_HH2_xy_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_resized_HH2_xy_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_resized_HH2_xy_blurred_In1_data : std_logic_vector(15 downto 0);
	signal ai_resized_HH2_xy_blurred_In1_send : std_logic;
	signal ai_resized_HH2_xy_blurred_In1_ack : std_logic;
	signal ai_resized_HH2_xy_blurred_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_resized_HH2_xy_blurred_Out1_data : std_logic_vector(15 downto 0);
	signal ao_resized_HH2_xy_blurred_Out1_send : std_logic;
	signal ao_resized_HH2_xy_blurred_Out1_ack : std_logic;
	signal ao_resized_HH2_xy_blurred_Out1_rdy : std_logic;
	signal ao_resized_HH2_xy_blurred_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_resized_HH2_xy_blurred_Out1_data : std_logic_vector(15 downto 0);
	signal aof_resized_HH2_xy_blurred_Out1_send : std_logic_vector(0 downto 0);
	signal aof_resized_HH2_xy_blurred_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_resized_HH2_xy_blurred_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_resized_HH2_xy_blurred_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_resized_HH3_xy_In1_data : std_logic_vector(15 downto 0);
	signal ai_resized_HH3_xy_In1_send : std_logic;
	signal ai_resized_HH3_xy_In1_ack : std_logic;
	signal ai_resized_HH3_xy_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_resized_HH3_xy_Out1_data : std_logic_vector(15 downto 0);
	signal ao_resized_HH3_xy_Out1_send : std_logic;
	signal ao_resized_HH3_xy_Out1_ack : std_logic;
	signal ao_resized_HH3_xy_Out1_rdy : std_logic;
	signal ao_resized_HH3_xy_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_resized_HH3_xy_Out1_data : std_logic_vector(15 downto 0);
	signal aof_resized_HH3_xy_Out1_send : std_logic_vector(0 downto 0);
	signal aof_resized_HH3_xy_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_resized_HH3_xy_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_resized_HH3_xy_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_resized_HH3_xy_blurred_In1_data : std_logic_vector(15 downto 0);
	signal ai_resized_HH3_xy_blurred_In1_send : std_logic;
	signal ai_resized_HH3_xy_blurred_In1_ack : std_logic;
	signal ai_resized_HH3_xy_blurred_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_resized_HH3_xy_blurred_Out1_data : std_logic_vector(15 downto 0);
	signal ao_resized_HH3_xy_blurred_Out1_send : std_logic;
	signal ao_resized_HH3_xy_blurred_Out1_ack : std_logic;
	signal ao_resized_HH3_xy_blurred_Out1_rdy : std_logic;
	signal ao_resized_HH3_xy_blurred_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_resized_HH3_xy_blurred_Out1_data : std_logic_vector(15 downto 0);
	signal aof_resized_HH3_xy_blurred_Out1_send : std_logic_vector(0 downto 0);
	signal aof_resized_HH3_xy_blurred_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_resized_HH3_xy_blurred_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_resized_HH3_xy_blurred_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_resized_LH1_xy_In1_data : std_logic_vector(15 downto 0);
	signal ai_resized_LH1_xy_In1_send : std_logic;
	signal ai_resized_LH1_xy_In1_ack : std_logic;
	signal ai_resized_LH1_xy_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_resized_LH1_xy_Out1_data : std_logic_vector(15 downto 0);
	signal ao_resized_LH1_xy_Out1_send : std_logic;
	signal ao_resized_LH1_xy_Out1_ack : std_logic;
	signal ao_resized_LH1_xy_Out1_rdy : std_logic;
	signal ao_resized_LH1_xy_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_resized_LH1_xy_Out1_data : std_logic_vector(15 downto 0);
	signal aof_resized_LH1_xy_Out1_send : std_logic_vector(0 downto 0);
	signal aof_resized_LH1_xy_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_resized_LH1_xy_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_resized_LH1_xy_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_resized_LH1_xy_blurred_In1_data : std_logic_vector(15 downto 0);
	signal ai_resized_LH1_xy_blurred_In1_send : std_logic;
	signal ai_resized_LH1_xy_blurred_In1_ack : std_logic;
	signal ai_resized_LH1_xy_blurred_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_resized_LH1_xy_blurred_Out1_data : std_logic_vector(15 downto 0);
	signal ao_resized_LH1_xy_blurred_Out1_send : std_logic;
	signal ao_resized_LH1_xy_blurred_Out1_ack : std_logic;
	signal ao_resized_LH1_xy_blurred_Out1_rdy : std_logic;
	signal ao_resized_LH1_xy_blurred_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_resized_LH1_xy_blurred_Out1_data : std_logic_vector(15 downto 0);
	signal aof_resized_LH1_xy_blurred_Out1_send : std_logic_vector(0 downto 0);
	signal aof_resized_LH1_xy_blurred_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_resized_LH1_xy_blurred_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_resized_LH1_xy_blurred_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_resized_LH2_xy_In1_data : std_logic_vector(15 downto 0);
	signal ai_resized_LH2_xy_In1_send : std_logic;
	signal ai_resized_LH2_xy_In1_ack : std_logic;
	signal ai_resized_LH2_xy_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_resized_LH2_xy_Out1_data : std_logic_vector(15 downto 0);
	signal ao_resized_LH2_xy_Out1_send : std_logic;
	signal ao_resized_LH2_xy_Out1_ack : std_logic;
	signal ao_resized_LH2_xy_Out1_rdy : std_logic;
	signal ao_resized_LH2_xy_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_resized_LH2_xy_Out1_data : std_logic_vector(15 downto 0);
	signal aof_resized_LH2_xy_Out1_send : std_logic_vector(0 downto 0);
	signal aof_resized_LH2_xy_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_resized_LH2_xy_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_resized_LH2_xy_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_resized_LH2_xy_blurred_In1_data : std_logic_vector(15 downto 0);
	signal ai_resized_LH2_xy_blurred_In1_send : std_logic;
	signal ai_resized_LH2_xy_blurred_In1_ack : std_logic;
	signal ai_resized_LH2_xy_blurred_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_resized_LH2_xy_blurred_Out1_data : std_logic_vector(15 downto 0);
	signal ao_resized_LH2_xy_blurred_Out1_send : std_logic;
	signal ao_resized_LH2_xy_blurred_Out1_ack : std_logic;
	signal ao_resized_LH2_xy_blurred_Out1_rdy : std_logic;
	signal ao_resized_LH2_xy_blurred_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_resized_LH2_xy_blurred_Out1_data : std_logic_vector(15 downto 0);
	signal aof_resized_LH2_xy_blurred_Out1_send : std_logic_vector(0 downto 0);
	signal aof_resized_LH2_xy_blurred_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_resized_LH2_xy_blurred_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_resized_LH2_xy_blurred_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_resized_LH3_xy_In1_data : std_logic_vector(15 downto 0);
	signal ai_resized_LH3_xy_In1_send : std_logic;
	signal ai_resized_LH3_xy_In1_ack : std_logic;
	signal ai_resized_LH3_xy_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_resized_LH3_xy_Out1_data : std_logic_vector(15 downto 0);
	signal ao_resized_LH3_xy_Out1_send : std_logic;
	signal ao_resized_LH3_xy_Out1_ack : std_logic;
	signal ao_resized_LH3_xy_Out1_rdy : std_logic;
	signal ao_resized_LH3_xy_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_resized_LH3_xy_Out1_data : std_logic_vector(15 downto 0);
	signal aof_resized_LH3_xy_Out1_send : std_logic_vector(0 downto 0);
	signal aof_resized_LH3_xy_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_resized_LH3_xy_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_resized_LH3_xy_Out1_count : std_logic_vector(15 downto 0);
	
	signal ai_resized_LH3_xy_blurred_In1_data : std_logic_vector(15 downto 0);
	signal ai_resized_LH3_xy_blurred_In1_send : std_logic;
	signal ai_resized_LH3_xy_blurred_In1_ack : std_logic;
	signal ai_resized_LH3_xy_blurred_In1_count : std_logic_vector(15 downto 0);
	
	signal ao_resized_LH3_xy_blurred_Out1_data : std_logic_vector(15 downto 0);
	signal ao_resized_LH3_xy_blurred_Out1_send : std_logic;
	signal ao_resized_LH3_xy_blurred_Out1_ack : std_logic;
	signal ao_resized_LH3_xy_blurred_Out1_rdy : std_logic;
	signal ao_resized_LH3_xy_blurred_Out1_count : std_logic_vector(15 downto 0);
	
	signal aof_resized_LH3_xy_blurred_Out1_data : std_logic_vector(15 downto 0);
	signal aof_resized_LH3_xy_blurred_Out1_send : std_logic_vector(0 downto 0);
	signal aof_resized_LH3_xy_blurred_Out1_ack : std_logic_vector(0 downto 0);
	signal aof_resized_LH3_xy_blurred_Out1_rdy : std_logic_vector(0 downto 0);
	signal aof_resized_LH3_xy_blurred_Out1_count : std_logic_vector(15 downto 0);

	-- --------------------------------------------------------------------------
	-- Network Instances
	-- --------------------------------------------------------------------------
	component LL1_H_iunzipFilter2D is
	port(
	     -- Instance LL1_H_iunzipFilter2D Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance LL1_H_iunzipFilter2D Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     Out2_data : out std_logic_vector(15 downto 0);
	     Out2_send : out std_logic;
	     Out2_ack : in std_logic;
	     Out2_rdy : in std_logic;
	     Out2_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component LL1_H_iunzipFilter2D;
	
	component HH1 is
	port(
	     -- Instance HH1 Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance HH1 Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component HH1;
	
	component LL2_H_iunzipFilter2D is
	port(
	     -- Instance LL2_H_iunzipFilter2D Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance LL2_H_iunzipFilter2D Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     Out2_data : out std_logic_vector(15 downto 0);
	     Out2_send : out std_logic;
	     Out2_ack : in std_logic;
	     Out2_rdy : in std_logic;
	     Out2_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component LL2_H_iunzipFilter2D;
	
	component HH2 is
	port(
	     -- Instance HH2 Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance HH2 Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component HH2;
	
	component LL3_H_iunzipFilter2D is
	port(
	     -- Instance LL3_H_iunzipFilter2D Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance LL3_H_iunzipFilter2D Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     Out2_data : out std_logic_vector(15 downto 0);
	     Out2_send : out std_logic;
	     Out2_ack : in std_logic;
	     Out2_rdy : in std_logic;
	     Out2_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component LL3_H_iunzipFilter2D;
	
	component HH3 is
	port(
	     -- Instance HH3 Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance HH3 Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component HH3;
	
	component HL1 is
	port(
	     -- Instance HL1 Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance HL1 Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component HL1;
	
	component HL2 is
	port(
	     -- Instance HL2 Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance HL2 Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component HL2;
	
	component HL3 is
	port(
	     -- Instance HL3 Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance HL3 Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component HL3;
	
	component LL1_L_iunzipFilter2D is
	port(
	     -- Instance LL1_L_iunzipFilter2D Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance LL1_L_iunzipFilter2D Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     Out2_data : out std_logic_vector(15 downto 0);
	     Out2_send : out std_logic;
	     Out2_ack : in std_logic;
	     Out2_rdy : in std_logic;
	     Out2_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component LL1_L_iunzipFilter2D;
	
	component LH1 is
	port(
	     -- Instance LH1 Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance LH1 Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component LH1;
	
	component LL2_L_iunzipFilter2D is
	port(
	     -- Instance LL2_L_iunzipFilter2D Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance LL2_L_iunzipFilter2D Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     Out2_data : out std_logic_vector(15 downto 0);
	     Out2_send : out std_logic;
	     Out2_ack : in std_logic;
	     Out2_rdy : in std_logic;
	     Out2_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component LL2_L_iunzipFilter2D;
	
	component LH2 is
	port(
	     -- Instance LH2 Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance LH2 Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component LH2;
	
	component LL3_L_iunzipFilter2D is
	port(
	     -- Instance LL3_L_iunzipFilter2D Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance LL3_L_iunzipFilter2D Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     Out2_data : out std_logic_vector(15 downto 0);
	     Out2_send : out std_logic;
	     Out2_ack : in std_logic;
	     Out2_rdy : in std_logic;
	     Out2_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component LL3_L_iunzipFilter2D;
	
	component LH3 is
	port(
	     -- Instance LH3 Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance LH3 Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component LH3;
	
	component LL1 is
	port(
	     -- Instance LL1 Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance LL1 Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component LL1;
	
	component image1_iunzip is
	port(
	     -- Instance image1_iunzip Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance image1_iunzip Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     Out2_data : out std_logic_vector(15 downto 0);
	     Out2_send : out std_logic;
	     Out2_ack : in std_logic;
	     Out2_rdy : in std_logic;
	     Out2_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component image1_iunzip;
	
	component LL1_H is
	port(
	     -- Instance LL1_H Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance LL1_H Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component LL1_H;
	
	component LL1_L is
	port(
	     -- Instance LL1_L Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance LL1_L Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component LL1_L;
	
	component LL2 is
	port(
	     -- Instance LL2 Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance LL2 Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component LL2;
	
	component LL1_iunzip is
	port(
	     -- Instance LL1_iunzip Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance LL1_iunzip Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     Out2_data : out std_logic_vector(15 downto 0);
	     Out2_send : out std_logic;
	     Out2_ack : in std_logic;
	     Out2_rdy : in std_logic;
	     Out2_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component LL1_iunzip;
	
	component LL2_H is
	port(
	     -- Instance LL2_H Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance LL2_H Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component LL2_H;
	
	component LL2_L is
	port(
	     -- Instance LL2_L Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance LL2_L Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component LL2_L;
	
	component LL3 is
	port(
	     -- Instance LL3 Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance LL3 Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component LL3;
	
	component LL2_iunzip is
	port(
	     -- Instance LL2_iunzip Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance LL2_iunzip Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     Out2_data : out std_logic_vector(15 downto 0);
	     Out2_send : out std_logic;
	     Out2_ack : in std_logic;
	     Out2_rdy : in std_logic;
	     Out2_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component LL2_iunzip;
	
	component LL3_H is
	port(
	     -- Instance LL3_H Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance LL3_H Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component LL3_H;
	
	component LL3_L is
	port(
	     -- Instance LL3_L Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance LL3_L Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component LL3_L;
	
	component image1 is
	port(
	     -- Instance image1 Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance image1 Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component image1;
	
	component mapDia is
	port(
	     -- Instance mapDia Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     In2_data : in std_logic_vector(15 downto 0);
	     In2_send : in std_logic;
	     In2_ack : out std_logic;
	     In2_count : in std_logic_vector(15 downto 0);
	     In3_data : in std_logic_vector(15 downto 0);
	     In3_send : in std_logic;
	     In3_ack : out std_logic;
	     In3_count : in std_logic_vector(15 downto 0);
	     -- Instance mapDia Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component mapDia;
	
	component mapFinal is
	port(
	     -- Instance mapFinal Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     In2_data : in std_logic_vector(15 downto 0);
	     In2_send : in std_logic;
	     In2_ack : out std_logic;
	     In2_count : in std_logic_vector(15 downto 0);
	     -- Instance mapFinal Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component mapFinal;
	
	component mapVer is
	port(
	     -- Instance mapVer Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     In2_data : in std_logic_vector(15 downto 0);
	     In2_send : in std_logic;
	     In2_ack : out std_logic;
	     In2_count : in std_logic_vector(15 downto 0);
	     In3_data : in std_logic_vector(15 downto 0);
	     In3_send : in std_logic;
	     In3_ack : out std_logic;
	     In3_count : in std_logic_vector(15 downto 0);
	     -- Instance mapVer Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component mapVer;
	
	component resized_HH1_xy is
	port(
	     -- Instance resized_HH1_xy Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance resized_HH1_xy Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component resized_HH1_xy;
	
	component resized_HH1_xy_blurred is
	port(
	     -- Instance resized_HH1_xy_blurred Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance resized_HH1_xy_blurred Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component resized_HH1_xy_blurred;
	
	component resized_HH2_xy is
	port(
	     -- Instance resized_HH2_xy Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance resized_HH2_xy Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component resized_HH2_xy;
	
	component resized_HH2_xy_blurred is
	port(
	     -- Instance resized_HH2_xy_blurred Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance resized_HH2_xy_blurred Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component resized_HH2_xy_blurred;
	
	component resized_HH3_xy is
	port(
	     -- Instance resized_HH3_xy Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance resized_HH3_xy Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component resized_HH3_xy;
	
	component resized_HH3_xy_blurred is
	port(
	     -- Instance resized_HH3_xy_blurred Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance resized_HH3_xy_blurred Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component resized_HH3_xy_blurred;
	
	component resized_LH1_xy is
	port(
	     -- Instance resized_LH1_xy Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance resized_LH1_xy Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component resized_LH1_xy;
	
	component resized_LH1_xy_blurred is
	port(
	     -- Instance resized_LH1_xy_blurred Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance resized_LH1_xy_blurred Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component resized_LH1_xy_blurred;
	
	component resized_LH2_xy is
	port(
	     -- Instance resized_LH2_xy Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance resized_LH2_xy Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component resized_LH2_xy;
	
	component resized_LH2_xy_blurred is
	port(
	     -- Instance resized_LH2_xy_blurred Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance resized_LH2_xy_blurred Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component resized_LH2_xy_blurred;
	
	component resized_LH3_xy is
	port(
	     -- Instance resized_LH3_xy Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance resized_LH3_xy Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component resized_LH3_xy;
	
	component resized_LH3_xy_blurred is
	port(
	     -- Instance resized_LH3_xy_blurred Input(s)
	     In1_data : in std_logic_vector(15 downto 0);
	     In1_send : in std_logic;
	     In1_ack : out std_logic;
	     In1_count : in std_logic_vector(15 downto 0);
	     -- Instance resized_LH3_xy_blurred Output(s)
	     Out1_data : out std_logic_vector(15 downto 0);
	     Out1_send : out std_logic;
	     Out1_ack : in std_logic;
	     Out1_rdy : in std_logic;
	     Out1_count : out std_logic_vector(15 downto 0);
	     clk: in std_logic;
	     reset: in std_logic);
	end component resized_LH3_xy_blurred;
	

begin
	-- Reset Controller
	rcon: entity SystemBuilder.resetController(behavioral)
	generic map(count => 1)
	port map( 
	         clocks => clocks, 
	         reset_in => reset, 
	         resets => resets);
	
	clocks(0) <= CLK;

	-- --------------------------------------------------------------------------
	-- Actor instances
	-- --------------------------------------------------------------------------
	i_LL1_H_iunzipFilter2D : component LL1_H_iunzipFilter2D
	port map(
		-- Instance LL1_H_iunzipFilter2D Input(s)
		In1_data => ai_LL1_H_iunzipFilter2D_In1_data,
		In1_send => ai_LL1_H_iunzipFilter2D_In1_send,
		In1_ack => ai_LL1_H_iunzipFilter2D_In1_ack,
		In1_count => ai_LL1_H_iunzipFilter2D_In1_count,
		-- Instance LL1_H_iunzipFilter2D Output(s)
		Out1_data => ao_LL1_H_iunzipFilter2D_Out1_data,
		Out1_send => ao_LL1_H_iunzipFilter2D_Out1_send,
		Out1_ack => ao_LL1_H_iunzipFilter2D_Out1_ack,
		Out1_rdy => ao_LL1_H_iunzipFilter2D_Out1_rdy,
		Out1_count => ao_LL1_H_iunzipFilter2D_Out1_count,
		
		Out2_data => ao_LL1_H_iunzipFilter2D_Out2_data,
		Out2_send => ao_LL1_H_iunzipFilter2D_Out2_send,
		Out2_ack => ao_LL1_H_iunzipFilter2D_Out2_ack,
		Out2_rdy => ao_LL1_H_iunzipFilter2D_Out2_rdy,
		Out2_count => ao_LL1_H_iunzipFilter2D_Out2_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_HH1 : component HH1
	port map(
		-- Instance HH1 Input(s)
		In1_data => ai_HH1_In1_data,
		In1_send => ai_HH1_In1_send,
		In1_ack => ai_HH1_In1_ack,
		In1_count => ai_HH1_In1_count,
		-- Instance HH1 Output(s)
		Out1_data => ao_HH1_Out1_data,
		Out1_send => ao_HH1_Out1_send,
		Out1_ack => ao_HH1_Out1_ack,
		Out1_rdy => ao_HH1_Out1_rdy,
		Out1_count => ao_HH1_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_LL2_H_iunzipFilter2D : component LL2_H_iunzipFilter2D
	port map(
		-- Instance LL2_H_iunzipFilter2D Input(s)
		In1_data => ai_LL2_H_iunzipFilter2D_In1_data,
		In1_send => ai_LL2_H_iunzipFilter2D_In1_send,
		In1_ack => ai_LL2_H_iunzipFilter2D_In1_ack,
		In1_count => ai_LL2_H_iunzipFilter2D_In1_count,
		-- Instance LL2_H_iunzipFilter2D Output(s)
		Out1_data => ao_LL2_H_iunzipFilter2D_Out1_data,
		Out1_send => ao_LL2_H_iunzipFilter2D_Out1_send,
		Out1_ack => ao_LL2_H_iunzipFilter2D_Out1_ack,
		Out1_rdy => ao_LL2_H_iunzipFilter2D_Out1_rdy,
		Out1_count => ao_LL2_H_iunzipFilter2D_Out1_count,
		
		Out2_data => ao_LL2_H_iunzipFilter2D_Out2_data,
		Out2_send => ao_LL2_H_iunzipFilter2D_Out2_send,
		Out2_ack => ao_LL2_H_iunzipFilter2D_Out2_ack,
		Out2_rdy => ao_LL2_H_iunzipFilter2D_Out2_rdy,
		Out2_count => ao_LL2_H_iunzipFilter2D_Out2_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_HH2 : component HH2
	port map(
		-- Instance HH2 Input(s)
		In1_data => ai_HH2_In1_data,
		In1_send => ai_HH2_In1_send,
		In1_ack => ai_HH2_In1_ack,
		In1_count => ai_HH2_In1_count,
		-- Instance HH2 Output(s)
		Out1_data => ao_HH2_Out1_data,
		Out1_send => ao_HH2_Out1_send,
		Out1_ack => ao_HH2_Out1_ack,
		Out1_rdy => ao_HH2_Out1_rdy,
		Out1_count => ao_HH2_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_LL3_H_iunzipFilter2D : component LL3_H_iunzipFilter2D
	port map(
		-- Instance LL3_H_iunzipFilter2D Input(s)
		In1_data => ai_LL3_H_iunzipFilter2D_In1_data,
		In1_send => ai_LL3_H_iunzipFilter2D_In1_send,
		In1_ack => ai_LL3_H_iunzipFilter2D_In1_ack,
		In1_count => ai_LL3_H_iunzipFilter2D_In1_count,
		-- Instance LL3_H_iunzipFilter2D Output(s)
		Out1_data => ao_LL3_H_iunzipFilter2D_Out1_data,
		Out1_send => ao_LL3_H_iunzipFilter2D_Out1_send,
		Out1_ack => ao_LL3_H_iunzipFilter2D_Out1_ack,
		Out1_rdy => ao_LL3_H_iunzipFilter2D_Out1_rdy,
		Out1_count => ao_LL3_H_iunzipFilter2D_Out1_count,
		
		Out2_data => ao_LL3_H_iunzipFilter2D_Out2_data,
		Out2_send => ao_LL3_H_iunzipFilter2D_Out2_send,
		Out2_ack => ao_LL3_H_iunzipFilter2D_Out2_ack,
		Out2_rdy => ao_LL3_H_iunzipFilter2D_Out2_rdy,
		Out2_count => ao_LL3_H_iunzipFilter2D_Out2_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_HH3 : component HH3
	port map(
		-- Instance HH3 Input(s)
		In1_data => ai_HH3_In1_data,
		In1_send => ai_HH3_In1_send,
		In1_ack => ai_HH3_In1_ack,
		In1_count => ai_HH3_In1_count,
		-- Instance HH3 Output(s)
		Out1_data => ao_HH3_Out1_data,
		Out1_send => ao_HH3_Out1_send,
		Out1_ack => ao_HH3_Out1_ack,
		Out1_rdy => ao_HH3_Out1_rdy,
		Out1_count => ao_HH3_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_HL1 : component HL1
	port map(
		-- Instance HL1 Input(s)
		In1_data => ai_HL1_In1_data,
		In1_send => ai_HL1_In1_send,
		In1_ack => ai_HL1_In1_ack,
		In1_count => ai_HL1_In1_count,
		-- Instance HL1 Output(s)
		Out1_data => ao_HL1_Out1_data,
		Out1_send => ao_HL1_Out1_send,
		Out1_ack => ao_HL1_Out1_ack,
		Out1_rdy => ao_HL1_Out1_rdy,
		Out1_count => ao_HL1_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_HL2 : component HL2
	port map(
		-- Instance HL2 Input(s)
		In1_data => ai_HL2_In1_data,
		In1_send => ai_HL2_In1_send,
		In1_ack => ai_HL2_In1_ack,
		In1_count => ai_HL2_In1_count,
		-- Instance HL2 Output(s)
		Out1_data => ao_HL2_Out1_data,
		Out1_send => ao_HL2_Out1_send,
		Out1_ack => ao_HL2_Out1_ack,
		Out1_rdy => ao_HL2_Out1_rdy,
		Out1_count => ao_HL2_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_HL3 : component HL3
	port map(
		-- Instance HL3 Input(s)
		In1_data => ai_HL3_In1_data,
		In1_send => ai_HL3_In1_send,
		In1_ack => ai_HL3_In1_ack,
		In1_count => ai_HL3_In1_count,
		-- Instance HL3 Output(s)
		Out1_data => ao_HL3_Out1_data,
		Out1_send => ao_HL3_Out1_send,
		Out1_ack => ao_HL3_Out1_ack,
		Out1_rdy => ao_HL3_Out1_rdy,
		Out1_count => ao_HL3_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_LL1_L_iunzipFilter2D : component LL1_L_iunzipFilter2D
	port map(
		-- Instance LL1_L_iunzipFilter2D Input(s)
		In1_data => ai_LL1_L_iunzipFilter2D_In1_data,
		In1_send => ai_LL1_L_iunzipFilter2D_In1_send,
		In1_ack => ai_LL1_L_iunzipFilter2D_In1_ack,
		In1_count => ai_LL1_L_iunzipFilter2D_In1_count,
		-- Instance LL1_L_iunzipFilter2D Output(s)
		Out1_data => ao_LL1_L_iunzipFilter2D_Out1_data,
		Out1_send => ao_LL1_L_iunzipFilter2D_Out1_send,
		Out1_ack => ao_LL1_L_iunzipFilter2D_Out1_ack,
		Out1_rdy => ao_LL1_L_iunzipFilter2D_Out1_rdy,
		Out1_count => ao_LL1_L_iunzipFilter2D_Out1_count,
		
		Out2_data => ao_LL1_L_iunzipFilter2D_Out2_data,
		Out2_send => ao_LL1_L_iunzipFilter2D_Out2_send,
		Out2_ack => ao_LL1_L_iunzipFilter2D_Out2_ack,
		Out2_rdy => ao_LL1_L_iunzipFilter2D_Out2_rdy,
		Out2_count => ao_LL1_L_iunzipFilter2D_Out2_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_LH1 : component LH1
	port map(
		-- Instance LH1 Input(s)
		In1_data => ai_LH1_In1_data,
		In1_send => ai_LH1_In1_send,
		In1_ack => ai_LH1_In1_ack,
		In1_count => ai_LH1_In1_count,
		-- Instance LH1 Output(s)
		Out1_data => ao_LH1_Out1_data,
		Out1_send => ao_LH1_Out1_send,
		Out1_ack => ao_LH1_Out1_ack,
		Out1_rdy => ao_LH1_Out1_rdy,
		Out1_count => ao_LH1_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_LL2_L_iunzipFilter2D : component LL2_L_iunzipFilter2D
	port map(
		-- Instance LL2_L_iunzipFilter2D Input(s)
		In1_data => ai_LL2_L_iunzipFilter2D_In1_data,
		In1_send => ai_LL2_L_iunzipFilter2D_In1_send,
		In1_ack => ai_LL2_L_iunzipFilter2D_In1_ack,
		In1_count => ai_LL2_L_iunzipFilter2D_In1_count,
		-- Instance LL2_L_iunzipFilter2D Output(s)
		Out1_data => ao_LL2_L_iunzipFilter2D_Out1_data,
		Out1_send => ao_LL2_L_iunzipFilter2D_Out1_send,
		Out1_ack => ao_LL2_L_iunzipFilter2D_Out1_ack,
		Out1_rdy => ao_LL2_L_iunzipFilter2D_Out1_rdy,
		Out1_count => ao_LL2_L_iunzipFilter2D_Out1_count,
		
		Out2_data => ao_LL2_L_iunzipFilter2D_Out2_data,
		Out2_send => ao_LL2_L_iunzipFilter2D_Out2_send,
		Out2_ack => ao_LL2_L_iunzipFilter2D_Out2_ack,
		Out2_rdy => ao_LL2_L_iunzipFilter2D_Out2_rdy,
		Out2_count => ao_LL2_L_iunzipFilter2D_Out2_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_LH2 : component LH2
	port map(
		-- Instance LH2 Input(s)
		In1_data => ai_LH2_In1_data,
		In1_send => ai_LH2_In1_send,
		In1_ack => ai_LH2_In1_ack,
		In1_count => ai_LH2_In1_count,
		-- Instance LH2 Output(s)
		Out1_data => ao_LH2_Out1_data,
		Out1_send => ao_LH2_Out1_send,
		Out1_ack => ao_LH2_Out1_ack,
		Out1_rdy => ao_LH2_Out1_rdy,
		Out1_count => ao_LH2_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_LL3_L_iunzipFilter2D : component LL3_L_iunzipFilter2D
	port map(
		-- Instance LL3_L_iunzipFilter2D Input(s)
		In1_data => ai_LL3_L_iunzipFilter2D_In1_data,
		In1_send => ai_LL3_L_iunzipFilter2D_In1_send,
		In1_ack => ai_LL3_L_iunzipFilter2D_In1_ack,
		In1_count => ai_LL3_L_iunzipFilter2D_In1_count,
		-- Instance LL3_L_iunzipFilter2D Output(s)
		Out1_data => ao_LL3_L_iunzipFilter2D_Out1_data,
		Out1_send => ao_LL3_L_iunzipFilter2D_Out1_send,
		Out1_ack => ao_LL3_L_iunzipFilter2D_Out1_ack,
		Out1_rdy => ao_LL3_L_iunzipFilter2D_Out1_rdy,
		Out1_count => ao_LL3_L_iunzipFilter2D_Out1_count,
		
		Out2_data => ao_LL3_L_iunzipFilter2D_Out2_data,
		Out2_send => ao_LL3_L_iunzipFilter2D_Out2_send,
		Out2_ack => ao_LL3_L_iunzipFilter2D_Out2_ack,
		Out2_rdy => ao_LL3_L_iunzipFilter2D_Out2_rdy,
		Out2_count => ao_LL3_L_iunzipFilter2D_Out2_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_LH3 : component LH3
	port map(
		-- Instance LH3 Input(s)
		In1_data => ai_LH3_In1_data,
		In1_send => ai_LH3_In1_send,
		In1_ack => ai_LH3_In1_ack,
		In1_count => ai_LH3_In1_count,
		-- Instance LH3 Output(s)
		Out1_data => ao_LH3_Out1_data,
		Out1_send => ao_LH3_Out1_send,
		Out1_ack => ao_LH3_Out1_ack,
		Out1_rdy => ao_LH3_Out1_rdy,
		Out1_count => ao_LH3_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_LL1 : component LL1
	port map(
		-- Instance LL1 Input(s)
		In1_data => ai_LL1_In1_data,
		In1_send => ai_LL1_In1_send,
		In1_ack => ai_LL1_In1_ack,
		In1_count => ai_LL1_In1_count,
		-- Instance LL1 Output(s)
		Out1_data => ao_LL1_Out1_data,
		Out1_send => ao_LL1_Out1_send,
		Out1_ack => ao_LL1_Out1_ack,
		Out1_rdy => ao_LL1_Out1_rdy,
		Out1_count => ao_LL1_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_image1_iunzip : component image1_iunzip
	port map(
		-- Instance image1_iunzip Input(s)
		In1_data => ai_image1_iunzip_In1_data,
		In1_send => ai_image1_iunzip_In1_send,
		In1_ack => ai_image1_iunzip_In1_ack,
		In1_count => ai_image1_iunzip_In1_count,
		-- Instance image1_iunzip Output(s)
		Out1_data => ao_image1_iunzip_Out1_data,
		Out1_send => ao_image1_iunzip_Out1_send,
		Out1_ack => ao_image1_iunzip_Out1_ack,
		Out1_rdy => ao_image1_iunzip_Out1_rdy,
		Out1_count => ao_image1_iunzip_Out1_count,
		
		Out2_data => ao_image1_iunzip_Out2_data,
		Out2_send => ao_image1_iunzip_Out2_send,
		Out2_ack => ao_image1_iunzip_Out2_ack,
		Out2_rdy => ao_image1_iunzip_Out2_rdy,
		Out2_count => ao_image1_iunzip_Out2_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_LL1_H : component LL1_H
	port map(
		-- Instance LL1_H Input(s)
		In1_data => ai_LL1_H_In1_data,
		In1_send => ai_LL1_H_In1_send,
		In1_ack => ai_LL1_H_In1_ack,
		In1_count => ai_LL1_H_In1_count,
		-- Instance LL1_H Output(s)
		Out1_data => ao_LL1_H_Out1_data,
		Out1_send => ao_LL1_H_Out1_send,
		Out1_ack => ao_LL1_H_Out1_ack,
		Out1_rdy => ao_LL1_H_Out1_rdy,
		Out1_count => ao_LL1_H_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_LL1_L : component LL1_L
	port map(
		-- Instance LL1_L Input(s)
		In1_data => ai_LL1_L_In1_data,
		In1_send => ai_LL1_L_In1_send,
		In1_ack => ai_LL1_L_In1_ack,
		In1_count => ai_LL1_L_In1_count,
		-- Instance LL1_L Output(s)
		Out1_data => ao_LL1_L_Out1_data,
		Out1_send => ao_LL1_L_Out1_send,
		Out1_ack => ao_LL1_L_Out1_ack,
		Out1_rdy => ao_LL1_L_Out1_rdy,
		Out1_count => ao_LL1_L_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_LL2 : component LL2
	port map(
		-- Instance LL2 Input(s)
		In1_data => ai_LL2_In1_data,
		In1_send => ai_LL2_In1_send,
		In1_ack => ai_LL2_In1_ack,
		In1_count => ai_LL2_In1_count,
		-- Instance LL2 Output(s)
		Out1_data => ao_LL2_Out1_data,
		Out1_send => ao_LL2_Out1_send,
		Out1_ack => ao_LL2_Out1_ack,
		Out1_rdy => ao_LL2_Out1_rdy,
		Out1_count => ao_LL2_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_LL1_iunzip : component LL1_iunzip
	port map(
		-- Instance LL1_iunzip Input(s)
		In1_data => ai_LL1_iunzip_In1_data,
		In1_send => ai_LL1_iunzip_In1_send,
		In1_ack => ai_LL1_iunzip_In1_ack,
		In1_count => ai_LL1_iunzip_In1_count,
		-- Instance LL1_iunzip Output(s)
		Out1_data => ao_LL1_iunzip_Out1_data,
		Out1_send => ao_LL1_iunzip_Out1_send,
		Out1_ack => ao_LL1_iunzip_Out1_ack,
		Out1_rdy => ao_LL1_iunzip_Out1_rdy,
		Out1_count => ao_LL1_iunzip_Out1_count,
		
		Out2_data => ao_LL1_iunzip_Out2_data,
		Out2_send => ao_LL1_iunzip_Out2_send,
		Out2_ack => ao_LL1_iunzip_Out2_ack,
		Out2_rdy => ao_LL1_iunzip_Out2_rdy,
		Out2_count => ao_LL1_iunzip_Out2_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_LL2_H : component LL2_H
	port map(
		-- Instance LL2_H Input(s)
		In1_data => ai_LL2_H_In1_data,
		In1_send => ai_LL2_H_In1_send,
		In1_ack => ai_LL2_H_In1_ack,
		In1_count => ai_LL2_H_In1_count,
		-- Instance LL2_H Output(s)
		Out1_data => ao_LL2_H_Out1_data,
		Out1_send => ao_LL2_H_Out1_send,
		Out1_ack => ao_LL2_H_Out1_ack,
		Out1_rdy => ao_LL2_H_Out1_rdy,
		Out1_count => ao_LL2_H_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_LL2_L : component LL2_L
	port map(
		-- Instance LL2_L Input(s)
		In1_data => ai_LL2_L_In1_data,
		In1_send => ai_LL2_L_In1_send,
		In1_ack => ai_LL2_L_In1_ack,
		In1_count => ai_LL2_L_In1_count,
		-- Instance LL2_L Output(s)
		Out1_data => ao_LL2_L_Out1_data,
		Out1_send => ao_LL2_L_Out1_send,
		Out1_ack => ao_LL2_L_Out1_ack,
		Out1_rdy => ao_LL2_L_Out1_rdy,
		Out1_count => ao_LL2_L_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_LL3 : component LL3
	port map(
		-- Instance LL3 Input(s)
		In1_data => ai_LL3_In1_data,
		In1_send => ai_LL3_In1_send,
		In1_ack => ai_LL3_In1_ack,
		In1_count => ai_LL3_In1_count,
		-- Instance LL3 Output(s)
		Out1_data => ao_LL3_Out1_data,
		Out1_send => ao_LL3_Out1_send,
		Out1_ack => ao_LL3_Out1_ack,
		Out1_rdy => ao_LL3_Out1_rdy,
		Out1_count => ao_LL3_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_LL2_iunzip : component LL2_iunzip
	port map(
		-- Instance LL2_iunzip Input(s)
		In1_data => ai_LL2_iunzip_In1_data,
		In1_send => ai_LL2_iunzip_In1_send,
		In1_ack => ai_LL2_iunzip_In1_ack,
		In1_count => ai_LL2_iunzip_In1_count,
		-- Instance LL2_iunzip Output(s)
		Out1_data => ao_LL2_iunzip_Out1_data,
		Out1_send => ao_LL2_iunzip_Out1_send,
		Out1_ack => ao_LL2_iunzip_Out1_ack,
		Out1_rdy => ao_LL2_iunzip_Out1_rdy,
		Out1_count => ao_LL2_iunzip_Out1_count,
		
		Out2_data => ao_LL2_iunzip_Out2_data,
		Out2_send => ao_LL2_iunzip_Out2_send,
		Out2_ack => ao_LL2_iunzip_Out2_ack,
		Out2_rdy => ao_LL2_iunzip_Out2_rdy,
		Out2_count => ao_LL2_iunzip_Out2_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_LL3_H : component LL3_H
	port map(
		-- Instance LL3_H Input(s)
		In1_data => ai_LL3_H_In1_data,
		In1_send => ai_LL3_H_In1_send,
		In1_ack => ai_LL3_H_In1_ack,
		In1_count => ai_LL3_H_In1_count,
		-- Instance LL3_H Output(s)
		Out1_data => ao_LL3_H_Out1_data,
		Out1_send => ao_LL3_H_Out1_send,
		Out1_ack => ao_LL3_H_Out1_ack,
		Out1_rdy => ao_LL3_H_Out1_rdy,
		Out1_count => ao_LL3_H_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_LL3_L : component LL3_L
	port map(
		-- Instance LL3_L Input(s)
		In1_data => ai_LL3_L_In1_data,
		In1_send => ai_LL3_L_In1_send,
		In1_ack => ai_LL3_L_In1_ack,
		In1_count => ai_LL3_L_In1_count,
		-- Instance LL3_L Output(s)
		Out1_data => ao_LL3_L_Out1_data,
		Out1_send => ao_LL3_L_Out1_send,
		Out1_ack => ao_LL3_L_Out1_ack,
		Out1_rdy => ao_LL3_L_Out1_rdy,
		Out1_count => ao_LL3_L_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_image1 : component image1
	port map(
		-- Instance image1 Input(s)
		In1_data => ai_image1_In1_data,
		In1_send => ai_image1_In1_send,
		In1_ack => ai_image1_In1_ack,
		In1_count => ai_image1_In1_count,
		-- Instance image1 Output(s)
		Out1_data => ao_image1_Out1_data,
		Out1_send => ao_image1_Out1_send,
		Out1_ack => ao_image1_Out1_ack,
		Out1_rdy => ao_image1_Out1_rdy,
		Out1_count => ao_image1_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_mapDia : component mapDia
	port map(
		-- Instance mapDia Input(s)
		In1_data => ai_mapDia_In1_data,
		In1_send => ai_mapDia_In1_send,
		In1_ack => ai_mapDia_In1_ack,
		In1_count => ai_mapDia_In1_count,
		
		In2_data => ai_mapDia_In2_data,
		In2_send => ai_mapDia_In2_send,
		In2_ack => ai_mapDia_In2_ack,
		In2_count => ai_mapDia_In2_count,
		
		In3_data => ai_mapDia_In3_data,
		In3_send => ai_mapDia_In3_send,
		In3_ack => ai_mapDia_In3_ack,
		In3_count => ai_mapDia_In3_count,
		-- Instance mapDia Output(s)
		Out1_data => ao_mapDia_Out1_data,
		Out1_send => ao_mapDia_Out1_send,
		Out1_ack => ao_mapDia_Out1_ack,
		Out1_rdy => ao_mapDia_Out1_rdy,
		Out1_count => ao_mapDia_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_mapFinal : component mapFinal
	port map(
		-- Instance mapFinal Input(s)
		In1_data => ai_mapFinal_In1_data,
		In1_send => ai_mapFinal_In1_send,
		In1_ack => ai_mapFinal_In1_ack,
		In1_count => ai_mapFinal_In1_count,
		
		In2_data => ai_mapFinal_In2_data,
		In2_send => ai_mapFinal_In2_send,
		In2_ack => ai_mapFinal_In2_ack,
		In2_count => ai_mapFinal_In2_count,
		-- Instance mapFinal Output(s)
		Out1_data => ao_mapFinal_Out1_data,
		Out1_send => ao_mapFinal_Out1_send,
		Out1_ack => ao_mapFinal_Out1_ack,
		Out1_rdy => ao_mapFinal_Out1_rdy,
		Out1_count => ao_mapFinal_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_mapVer : component mapVer
	port map(
		-- Instance mapVer Input(s)
		In1_data => ai_mapVer_In1_data,
		In1_send => ai_mapVer_In1_send,
		In1_ack => ai_mapVer_In1_ack,
		In1_count => ai_mapVer_In1_count,
		
		In2_data => ai_mapVer_In2_data,
		In2_send => ai_mapVer_In2_send,
		In2_ack => ai_mapVer_In2_ack,
		In2_count => ai_mapVer_In2_count,
		
		In3_data => ai_mapVer_In3_data,
		In3_send => ai_mapVer_In3_send,
		In3_ack => ai_mapVer_In3_ack,
		In3_count => ai_mapVer_In3_count,
		-- Instance mapVer Output(s)
		Out1_data => ao_mapVer_Out1_data,
		Out1_send => ao_mapVer_Out1_send,
		Out1_ack => ao_mapVer_Out1_ack,
		Out1_rdy => ao_mapVer_Out1_rdy,
		Out1_count => ao_mapVer_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_resized_HH1_xy : component resized_HH1_xy
	port map(
		-- Instance resized_HH1_xy Input(s)
		In1_data => ai_resized_HH1_xy_In1_data,
		In1_send => ai_resized_HH1_xy_In1_send,
		In1_ack => ai_resized_HH1_xy_In1_ack,
		In1_count => ai_resized_HH1_xy_In1_count,
		-- Instance resized_HH1_xy Output(s)
		Out1_data => ao_resized_HH1_xy_Out1_data,
		Out1_send => ao_resized_HH1_xy_Out1_send,
		Out1_ack => ao_resized_HH1_xy_Out1_ack,
		Out1_rdy => ao_resized_HH1_xy_Out1_rdy,
		Out1_count => ao_resized_HH1_xy_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_resized_HH1_xy_blurred : component resized_HH1_xy_blurred
	port map(
		-- Instance resized_HH1_xy_blurred Input(s)
		In1_data => ai_resized_HH1_xy_blurred_In1_data,
		In1_send => ai_resized_HH1_xy_blurred_In1_send,
		In1_ack => ai_resized_HH1_xy_blurred_In1_ack,
		In1_count => ai_resized_HH1_xy_blurred_In1_count,
		-- Instance resized_HH1_xy_blurred Output(s)
		Out1_data => ao_resized_HH1_xy_blurred_Out1_data,
		Out1_send => ao_resized_HH1_xy_blurred_Out1_send,
		Out1_ack => ao_resized_HH1_xy_blurred_Out1_ack,
		Out1_rdy => ao_resized_HH1_xy_blurred_Out1_rdy,
		Out1_count => ao_resized_HH1_xy_blurred_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_resized_HH2_xy : component resized_HH2_xy
	port map(
		-- Instance resized_HH2_xy Input(s)
		In1_data => ai_resized_HH2_xy_In1_data,
		In1_send => ai_resized_HH2_xy_In1_send,
		In1_ack => ai_resized_HH2_xy_In1_ack,
		In1_count => ai_resized_HH2_xy_In1_count,
		-- Instance resized_HH2_xy Output(s)
		Out1_data => ao_resized_HH2_xy_Out1_data,
		Out1_send => ao_resized_HH2_xy_Out1_send,
		Out1_ack => ao_resized_HH2_xy_Out1_ack,
		Out1_rdy => ao_resized_HH2_xy_Out1_rdy,
		Out1_count => ao_resized_HH2_xy_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_resized_HH2_xy_blurred : component resized_HH2_xy_blurred
	port map(
		-- Instance resized_HH2_xy_blurred Input(s)
		In1_data => ai_resized_HH2_xy_blurred_In1_data,
		In1_send => ai_resized_HH2_xy_blurred_In1_send,
		In1_ack => ai_resized_HH2_xy_blurred_In1_ack,
		In1_count => ai_resized_HH2_xy_blurred_In1_count,
		-- Instance resized_HH2_xy_blurred Output(s)
		Out1_data => ao_resized_HH2_xy_blurred_Out1_data,
		Out1_send => ao_resized_HH2_xy_blurred_Out1_send,
		Out1_ack => ao_resized_HH2_xy_blurred_Out1_ack,
		Out1_rdy => ao_resized_HH2_xy_blurred_Out1_rdy,
		Out1_count => ao_resized_HH2_xy_blurred_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_resized_HH3_xy : component resized_HH3_xy
	port map(
		-- Instance resized_HH3_xy Input(s)
		In1_data => ai_resized_HH3_xy_In1_data,
		In1_send => ai_resized_HH3_xy_In1_send,
		In1_ack => ai_resized_HH3_xy_In1_ack,
		In1_count => ai_resized_HH3_xy_In1_count,
		-- Instance resized_HH3_xy Output(s)
		Out1_data => ao_resized_HH3_xy_Out1_data,
		Out1_send => ao_resized_HH3_xy_Out1_send,
		Out1_ack => ao_resized_HH3_xy_Out1_ack,
		Out1_rdy => ao_resized_HH3_xy_Out1_rdy,
		Out1_count => ao_resized_HH3_xy_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_resized_HH3_xy_blurred : component resized_HH3_xy_blurred
	port map(
		-- Instance resized_HH3_xy_blurred Input(s)
		In1_data => ai_resized_HH3_xy_blurred_In1_data,
		In1_send => ai_resized_HH3_xy_blurred_In1_send,
		In1_ack => ai_resized_HH3_xy_blurred_In1_ack,
		In1_count => ai_resized_HH3_xy_blurred_In1_count,
		-- Instance resized_HH3_xy_blurred Output(s)
		Out1_data => ao_resized_HH3_xy_blurred_Out1_data,
		Out1_send => ao_resized_HH3_xy_blurred_Out1_send,
		Out1_ack => ao_resized_HH3_xy_blurred_Out1_ack,
		Out1_rdy => ao_resized_HH3_xy_blurred_Out1_rdy,
		Out1_count => ao_resized_HH3_xy_blurred_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_resized_LH1_xy : component resized_LH1_xy
	port map(
		-- Instance resized_LH1_xy Input(s)
		In1_data => ai_resized_LH1_xy_In1_data,
		In1_send => ai_resized_LH1_xy_In1_send,
		In1_ack => ai_resized_LH1_xy_In1_ack,
		In1_count => ai_resized_LH1_xy_In1_count,
		-- Instance resized_LH1_xy Output(s)
		Out1_data => ao_resized_LH1_xy_Out1_data,
		Out1_send => ao_resized_LH1_xy_Out1_send,
		Out1_ack => ao_resized_LH1_xy_Out1_ack,
		Out1_rdy => ao_resized_LH1_xy_Out1_rdy,
		Out1_count => ao_resized_LH1_xy_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_resized_LH1_xy_blurred : component resized_LH1_xy_blurred
	port map(
		-- Instance resized_LH1_xy_blurred Input(s)
		In1_data => ai_resized_LH1_xy_blurred_In1_data,
		In1_send => ai_resized_LH1_xy_blurred_In1_send,
		In1_ack => ai_resized_LH1_xy_blurred_In1_ack,
		In1_count => ai_resized_LH1_xy_blurred_In1_count,
		-- Instance resized_LH1_xy_blurred Output(s)
		Out1_data => ao_resized_LH1_xy_blurred_Out1_data,
		Out1_send => ao_resized_LH1_xy_blurred_Out1_send,
		Out1_ack => ao_resized_LH1_xy_blurred_Out1_ack,
		Out1_rdy => ao_resized_LH1_xy_blurred_Out1_rdy,
		Out1_count => ao_resized_LH1_xy_blurred_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_resized_LH2_xy : component resized_LH2_xy
	port map(
		-- Instance resized_LH2_xy Input(s)
		In1_data => ai_resized_LH2_xy_In1_data,
		In1_send => ai_resized_LH2_xy_In1_send,
		In1_ack => ai_resized_LH2_xy_In1_ack,
		In1_count => ai_resized_LH2_xy_In1_count,
		-- Instance resized_LH2_xy Output(s)
		Out1_data => ao_resized_LH2_xy_Out1_data,
		Out1_send => ao_resized_LH2_xy_Out1_send,
		Out1_ack => ao_resized_LH2_xy_Out1_ack,
		Out1_rdy => ao_resized_LH2_xy_Out1_rdy,
		Out1_count => ao_resized_LH2_xy_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_resized_LH2_xy_blurred : component resized_LH2_xy_blurred
	port map(
		-- Instance resized_LH2_xy_blurred Input(s)
		In1_data => ai_resized_LH2_xy_blurred_In1_data,
		In1_send => ai_resized_LH2_xy_blurred_In1_send,
		In1_ack => ai_resized_LH2_xy_blurred_In1_ack,
		In1_count => ai_resized_LH2_xy_blurred_In1_count,
		-- Instance resized_LH2_xy_blurred Output(s)
		Out1_data => ao_resized_LH2_xy_blurred_Out1_data,
		Out1_send => ao_resized_LH2_xy_blurred_Out1_send,
		Out1_ack => ao_resized_LH2_xy_blurred_Out1_ack,
		Out1_rdy => ao_resized_LH2_xy_blurred_Out1_rdy,
		Out1_count => ao_resized_LH2_xy_blurred_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_resized_LH3_xy : component resized_LH3_xy
	port map(
		-- Instance resized_LH3_xy Input(s)
		In1_data => ai_resized_LH3_xy_In1_data,
		In1_send => ai_resized_LH3_xy_In1_send,
		In1_ack => ai_resized_LH3_xy_In1_ack,
		In1_count => ai_resized_LH3_xy_In1_count,
		-- Instance resized_LH3_xy Output(s)
		Out1_data => ao_resized_LH3_xy_Out1_data,
		Out1_send => ao_resized_LH3_xy_Out1_send,
		Out1_ack => ao_resized_LH3_xy_Out1_ack,
		Out1_rdy => ao_resized_LH3_xy_Out1_rdy,
		Out1_count => ao_resized_LH3_xy_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	i_resized_LH3_xy_blurred : component resized_LH3_xy_blurred
	port map(
		-- Instance resized_LH3_xy_blurred Input(s)
		In1_data => ai_resized_LH3_xy_blurred_In1_data,
		In1_send => ai_resized_LH3_xy_blurred_In1_send,
		In1_ack => ai_resized_LH3_xy_blurred_In1_ack,
		In1_count => ai_resized_LH3_xy_blurred_In1_count,
		-- Instance resized_LH3_xy_blurred Output(s)
		Out1_data => ao_resized_LH3_xy_blurred_Out1_data,
		Out1_send => ao_resized_LH3_xy_blurred_Out1_send,
		Out1_ack => ao_resized_LH3_xy_blurred_Out1_ack,
		Out1_rdy => ao_resized_LH3_xy_blurred_Out1_rdy,
		Out1_count => ao_resized_LH3_xy_blurred_Out1_count,
		-- Clock and Reset
	clk => clocks(0),
	--clk => clocks(0),
	reset => resets(0));
	
	-- --------------------------------------------------------------------------
	-- Nework Input Fanouts
	-- --------------------------------------------------------------------------
	f_ni_In : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ni_In_data,
		In_send => ni_In_send,
		In_ack => ni_In_ack,
		In_rdy => ni_In_rdy,
		In_count => ni_In_count,
		-- Fanout Out
		Out_data => nif_In_data,
		Out_send => nif_In_send,
		Out_ack => nif_In_ack,
		Out_rdy => nif_In_rdy,
		Out_count => nif_In_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));

	-- --------------------------------------------------------------------------
	-- Actor Output Fanouts
	-- --------------------------------------------------------------------------
	f_ao_LL1_H_iunzipFilter2D_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_LL1_H_iunzipFilter2D_Out1_data,
		In_send => ao_LL1_H_iunzipFilter2D_Out1_send,
		In_ack => ao_LL1_H_iunzipFilter2D_Out1_ack,
		In_rdy => ao_LL1_H_iunzipFilter2D_Out1_rdy,
		In_count => ao_LL1_H_iunzipFilter2D_Out1_count,
		-- Fanout Out
		Out_data => aof_LL1_H_iunzipFilter2D_Out1_data,
		Out_send => aof_LL1_H_iunzipFilter2D_Out1_send,
		Out_ack => aof_LL1_H_iunzipFilter2D_Out1_ack,
		Out_rdy => aof_LL1_H_iunzipFilter2D_Out1_rdy,
		Out_count => aof_LL1_H_iunzipFilter2D_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	f_ao_LL1_H_iunzipFilter2D_Out2 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_LL1_H_iunzipFilter2D_Out2_data,
		In_send => ao_LL1_H_iunzipFilter2D_Out2_send,
		In_ack => ao_LL1_H_iunzipFilter2D_Out2_ack,
		In_rdy => ao_LL1_H_iunzipFilter2D_Out2_rdy,
		In_count => ao_LL1_H_iunzipFilter2D_Out2_count,
		-- Fanout Out
		Out_data => aof_LL1_H_iunzipFilter2D_Out2_data,
		Out_send => aof_LL1_H_iunzipFilter2D_Out2_send,
		Out_ack => aof_LL1_H_iunzipFilter2D_Out2_ack,
		Out_rdy => aof_LL1_H_iunzipFilter2D_Out2_rdy,
		Out_count => aof_LL1_H_iunzipFilter2D_Out2_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_HH1_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_HH1_Out1_data,
		In_send => ao_HH1_Out1_send,
		In_ack => ao_HH1_Out1_ack,
		In_rdy => ao_HH1_Out1_rdy,
		In_count => ao_HH1_Out1_count,
		-- Fanout Out
		Out_data => aof_HH1_Out1_data,
		Out_send => aof_HH1_Out1_send,
		Out_ack => aof_HH1_Out1_ack,
		Out_rdy => aof_HH1_Out1_rdy,
		Out_count => aof_HH1_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_LL2_H_iunzipFilter2D_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_LL2_H_iunzipFilter2D_Out1_data,
		In_send => ao_LL2_H_iunzipFilter2D_Out1_send,
		In_ack => ao_LL2_H_iunzipFilter2D_Out1_ack,
		In_rdy => ao_LL2_H_iunzipFilter2D_Out1_rdy,
		In_count => ao_LL2_H_iunzipFilter2D_Out1_count,
		-- Fanout Out
		Out_data => aof_LL2_H_iunzipFilter2D_Out1_data,
		Out_send => aof_LL2_H_iunzipFilter2D_Out1_send,
		Out_ack => aof_LL2_H_iunzipFilter2D_Out1_ack,
		Out_rdy => aof_LL2_H_iunzipFilter2D_Out1_rdy,
		Out_count => aof_LL2_H_iunzipFilter2D_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	f_ao_LL2_H_iunzipFilter2D_Out2 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_LL2_H_iunzipFilter2D_Out2_data,
		In_send => ao_LL2_H_iunzipFilter2D_Out2_send,
		In_ack => ao_LL2_H_iunzipFilter2D_Out2_ack,
		In_rdy => ao_LL2_H_iunzipFilter2D_Out2_rdy,
		In_count => ao_LL2_H_iunzipFilter2D_Out2_count,
		-- Fanout Out
		Out_data => aof_LL2_H_iunzipFilter2D_Out2_data,
		Out_send => aof_LL2_H_iunzipFilter2D_Out2_send,
		Out_ack => aof_LL2_H_iunzipFilter2D_Out2_ack,
		Out_rdy => aof_LL2_H_iunzipFilter2D_Out2_rdy,
		Out_count => aof_LL2_H_iunzipFilter2D_Out2_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_HH2_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_HH2_Out1_data,
		In_send => ao_HH2_Out1_send,
		In_ack => ao_HH2_Out1_ack,
		In_rdy => ao_HH2_Out1_rdy,
		In_count => ao_HH2_Out1_count,
		-- Fanout Out
		Out_data => aof_HH2_Out1_data,
		Out_send => aof_HH2_Out1_send,
		Out_ack => aof_HH2_Out1_ack,
		Out_rdy => aof_HH2_Out1_rdy,
		Out_count => aof_HH2_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_LL3_H_iunzipFilter2D_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_LL3_H_iunzipFilter2D_Out1_data,
		In_send => ao_LL3_H_iunzipFilter2D_Out1_send,
		In_ack => ao_LL3_H_iunzipFilter2D_Out1_ack,
		In_rdy => ao_LL3_H_iunzipFilter2D_Out1_rdy,
		In_count => ao_LL3_H_iunzipFilter2D_Out1_count,
		-- Fanout Out
		Out_data => aof_LL3_H_iunzipFilter2D_Out1_data,
		Out_send => aof_LL3_H_iunzipFilter2D_Out1_send,
		Out_ack => aof_LL3_H_iunzipFilter2D_Out1_ack,
		Out_rdy => aof_LL3_H_iunzipFilter2D_Out1_rdy,
		Out_count => aof_LL3_H_iunzipFilter2D_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	f_ao_LL3_H_iunzipFilter2D_Out2 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_LL3_H_iunzipFilter2D_Out2_data,
		In_send => ao_LL3_H_iunzipFilter2D_Out2_send,
		In_ack => ao_LL3_H_iunzipFilter2D_Out2_ack,
		In_rdy => ao_LL3_H_iunzipFilter2D_Out2_rdy,
		In_count => ao_LL3_H_iunzipFilter2D_Out2_count,
		-- Fanout Out
		Out_data => aof_LL3_H_iunzipFilter2D_Out2_data,
		Out_send => aof_LL3_H_iunzipFilter2D_Out2_send,
		Out_ack => aof_LL3_H_iunzipFilter2D_Out2_ack,
		Out_rdy => aof_LL3_H_iunzipFilter2D_Out2_rdy,
		Out_count => aof_LL3_H_iunzipFilter2D_Out2_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_HH3_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_HH3_Out1_data,
		In_send => ao_HH3_Out1_send,
		In_ack => ao_HH3_Out1_ack,
		In_rdy => ao_HH3_Out1_rdy,
		In_count => ao_HH3_Out1_count,
		-- Fanout Out
		Out_data => aof_HH3_Out1_data,
		Out_send => aof_HH3_Out1_send,
		Out_ack => aof_HH3_Out1_ack,
		Out_rdy => aof_HH3_Out1_rdy,
		Out_count => aof_HH3_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_HL1_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_HL1_Out1_data,
		In_send => ao_HL1_Out1_send,
		In_ack => ao_HL1_Out1_ack,
		In_rdy => ao_HL1_Out1_rdy,
		In_count => ao_HL1_Out1_count,
		-- Fanout Out
		Out_data => aof_HL1_Out1_data,
		Out_send => aof_HL1_Out1_send,
		Out_ack => aof_HL1_Out1_ack,
		Out_rdy => aof_HL1_Out1_rdy,
		Out_count => aof_HL1_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_HL2_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_HL2_Out1_data,
		In_send => ao_HL2_Out1_send,
		In_ack => ao_HL2_Out1_ack,
		In_rdy => ao_HL2_Out1_rdy,
		In_count => ao_HL2_Out1_count,
		-- Fanout Out
		Out_data => aof_HL2_Out1_data,
		Out_send => aof_HL2_Out1_send,
		Out_ack => aof_HL2_Out1_ack,
		Out_rdy => aof_HL2_Out1_rdy,
		Out_count => aof_HL2_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_HL3_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_HL3_Out1_data,
		In_send => ao_HL3_Out1_send,
		In_ack => ao_HL3_Out1_ack,
		In_rdy => ao_HL3_Out1_rdy,
		In_count => ao_HL3_Out1_count,
		-- Fanout Out
		Out_data => aof_HL3_Out1_data,
		Out_send => aof_HL3_Out1_send,
		Out_ack => aof_HL3_Out1_ack,
		Out_rdy => aof_HL3_Out1_rdy,
		Out_count => aof_HL3_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_LL1_L_iunzipFilter2D_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_LL1_L_iunzipFilter2D_Out1_data,
		In_send => ao_LL1_L_iunzipFilter2D_Out1_send,
		In_ack => ao_LL1_L_iunzipFilter2D_Out1_ack,
		In_rdy => ao_LL1_L_iunzipFilter2D_Out1_rdy,
		In_count => ao_LL1_L_iunzipFilter2D_Out1_count,
		-- Fanout Out
		Out_data => aof_LL1_L_iunzipFilter2D_Out1_data,
		Out_send => aof_LL1_L_iunzipFilter2D_Out1_send,
		Out_ack => aof_LL1_L_iunzipFilter2D_Out1_ack,
		Out_rdy => aof_LL1_L_iunzipFilter2D_Out1_rdy,
		Out_count => aof_LL1_L_iunzipFilter2D_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	f_ao_LL1_L_iunzipFilter2D_Out2 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_LL1_L_iunzipFilter2D_Out2_data,
		In_send => ao_LL1_L_iunzipFilter2D_Out2_send,
		In_ack => ao_LL1_L_iunzipFilter2D_Out2_ack,
		In_rdy => ao_LL1_L_iunzipFilter2D_Out2_rdy,
		In_count => ao_LL1_L_iunzipFilter2D_Out2_count,
		-- Fanout Out
		Out_data => aof_LL1_L_iunzipFilter2D_Out2_data,
		Out_send => aof_LL1_L_iunzipFilter2D_Out2_send,
		Out_ack => aof_LL1_L_iunzipFilter2D_Out2_ack,
		Out_rdy => aof_LL1_L_iunzipFilter2D_Out2_rdy,
		Out_count => aof_LL1_L_iunzipFilter2D_Out2_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_LH1_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_LH1_Out1_data,
		In_send => ao_LH1_Out1_send,
		In_ack => ao_LH1_Out1_ack,
		In_rdy => ao_LH1_Out1_rdy,
		In_count => ao_LH1_Out1_count,
		-- Fanout Out
		Out_data => aof_LH1_Out1_data,
		Out_send => aof_LH1_Out1_send,
		Out_ack => aof_LH1_Out1_ack,
		Out_rdy => aof_LH1_Out1_rdy,
		Out_count => aof_LH1_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_LL2_L_iunzipFilter2D_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_LL2_L_iunzipFilter2D_Out1_data,
		In_send => ao_LL2_L_iunzipFilter2D_Out1_send,
		In_ack => ao_LL2_L_iunzipFilter2D_Out1_ack,
		In_rdy => ao_LL2_L_iunzipFilter2D_Out1_rdy,
		In_count => ao_LL2_L_iunzipFilter2D_Out1_count,
		-- Fanout Out
		Out_data => aof_LL2_L_iunzipFilter2D_Out1_data,
		Out_send => aof_LL2_L_iunzipFilter2D_Out1_send,
		Out_ack => aof_LL2_L_iunzipFilter2D_Out1_ack,
		Out_rdy => aof_LL2_L_iunzipFilter2D_Out1_rdy,
		Out_count => aof_LL2_L_iunzipFilter2D_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	f_ao_LL2_L_iunzipFilter2D_Out2 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_LL2_L_iunzipFilter2D_Out2_data,
		In_send => ao_LL2_L_iunzipFilter2D_Out2_send,
		In_ack => ao_LL2_L_iunzipFilter2D_Out2_ack,
		In_rdy => ao_LL2_L_iunzipFilter2D_Out2_rdy,
		In_count => ao_LL2_L_iunzipFilter2D_Out2_count,
		-- Fanout Out
		Out_data => aof_LL2_L_iunzipFilter2D_Out2_data,
		Out_send => aof_LL2_L_iunzipFilter2D_Out2_send,
		Out_ack => aof_LL2_L_iunzipFilter2D_Out2_ack,
		Out_rdy => aof_LL2_L_iunzipFilter2D_Out2_rdy,
		Out_count => aof_LL2_L_iunzipFilter2D_Out2_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_LH2_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_LH2_Out1_data,
		In_send => ao_LH2_Out1_send,
		In_ack => ao_LH2_Out1_ack,
		In_rdy => ao_LH2_Out1_rdy,
		In_count => ao_LH2_Out1_count,
		-- Fanout Out
		Out_data => aof_LH2_Out1_data,
		Out_send => aof_LH2_Out1_send,
		Out_ack => aof_LH2_Out1_ack,
		Out_rdy => aof_LH2_Out1_rdy,
		Out_count => aof_LH2_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_LL3_L_iunzipFilter2D_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_LL3_L_iunzipFilter2D_Out1_data,
		In_send => ao_LL3_L_iunzipFilter2D_Out1_send,
		In_ack => ao_LL3_L_iunzipFilter2D_Out1_ack,
		In_rdy => ao_LL3_L_iunzipFilter2D_Out1_rdy,
		In_count => ao_LL3_L_iunzipFilter2D_Out1_count,
		-- Fanout Out
		Out_data => aof_LL3_L_iunzipFilter2D_Out1_data,
		Out_send => aof_LL3_L_iunzipFilter2D_Out1_send,
		Out_ack => aof_LL3_L_iunzipFilter2D_Out1_ack,
		Out_rdy => aof_LL3_L_iunzipFilter2D_Out1_rdy,
		Out_count => aof_LL3_L_iunzipFilter2D_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	f_ao_LL3_L_iunzipFilter2D_Out2 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_LL3_L_iunzipFilter2D_Out2_data,
		In_send => ao_LL3_L_iunzipFilter2D_Out2_send,
		In_ack => ao_LL3_L_iunzipFilter2D_Out2_ack,
		In_rdy => ao_LL3_L_iunzipFilter2D_Out2_rdy,
		In_count => ao_LL3_L_iunzipFilter2D_Out2_count,
		-- Fanout Out
		Out_data => aof_LL3_L_iunzipFilter2D_Out2_data,
		Out_send => aof_LL3_L_iunzipFilter2D_Out2_send,
		Out_ack => aof_LL3_L_iunzipFilter2D_Out2_ack,
		Out_rdy => aof_LL3_L_iunzipFilter2D_Out2_rdy,
		Out_count => aof_LL3_L_iunzipFilter2D_Out2_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_LH3_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_LH3_Out1_data,
		In_send => ao_LH3_Out1_send,
		In_ack => ao_LH3_Out1_ack,
		In_rdy => ao_LH3_Out1_rdy,
		In_count => ao_LH3_Out1_count,
		-- Fanout Out
		Out_data => aof_LH3_Out1_data,
		Out_send => aof_LH3_Out1_send,
		Out_ack => aof_LH3_Out1_ack,
		Out_rdy => aof_LH3_Out1_rdy,
		Out_count => aof_LH3_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_LL1_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_LL1_Out1_data,
		In_send => ao_LL1_Out1_send,
		In_ack => ao_LL1_Out1_ack,
		In_rdy => ao_LL1_Out1_rdy,
		In_count => ao_LL1_Out1_count,
		-- Fanout Out
		Out_data => aof_LL1_Out1_data,
		Out_send => aof_LL1_Out1_send,
		Out_ack => aof_LL1_Out1_ack,
		Out_rdy => aof_LL1_Out1_rdy,
		Out_count => aof_LL1_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_image1_iunzip_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_image1_iunzip_Out1_data,
		In_send => ao_image1_iunzip_Out1_send,
		In_ack => ao_image1_iunzip_Out1_ack,
		In_rdy => ao_image1_iunzip_Out1_rdy,
		In_count => ao_image1_iunzip_Out1_count,
		-- Fanout Out
		Out_data => aof_image1_iunzip_Out1_data,
		Out_send => aof_image1_iunzip_Out1_send,
		Out_ack => aof_image1_iunzip_Out1_ack,
		Out_rdy => aof_image1_iunzip_Out1_rdy,
		Out_count => aof_image1_iunzip_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	f_ao_image1_iunzip_Out2 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_image1_iunzip_Out2_data,
		In_send => ao_image1_iunzip_Out2_send,
		In_ack => ao_image1_iunzip_Out2_ack,
		In_rdy => ao_image1_iunzip_Out2_rdy,
		In_count => ao_image1_iunzip_Out2_count,
		-- Fanout Out
		Out_data => aof_image1_iunzip_Out2_data,
		Out_send => aof_image1_iunzip_Out2_send,
		Out_ack => aof_image1_iunzip_Out2_ack,
		Out_rdy => aof_image1_iunzip_Out2_rdy,
		Out_count => aof_image1_iunzip_Out2_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_LL1_H_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_LL1_H_Out1_data,
		In_send => ao_LL1_H_Out1_send,
		In_ack => ao_LL1_H_Out1_ack,
		In_rdy => ao_LL1_H_Out1_rdy,
		In_count => ao_LL1_H_Out1_count,
		-- Fanout Out
		Out_data => aof_LL1_H_Out1_data,
		Out_send => aof_LL1_H_Out1_send,
		Out_ack => aof_LL1_H_Out1_ack,
		Out_rdy => aof_LL1_H_Out1_rdy,
		Out_count => aof_LL1_H_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_LL1_L_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_LL1_L_Out1_data,
		In_send => ao_LL1_L_Out1_send,
		In_ack => ao_LL1_L_Out1_ack,
		In_rdy => ao_LL1_L_Out1_rdy,
		In_count => ao_LL1_L_Out1_count,
		-- Fanout Out
		Out_data => aof_LL1_L_Out1_data,
		Out_send => aof_LL1_L_Out1_send,
		Out_ack => aof_LL1_L_Out1_ack,
		Out_rdy => aof_LL1_L_Out1_rdy,
		Out_count => aof_LL1_L_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_LL2_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_LL2_Out1_data,
		In_send => ao_LL2_Out1_send,
		In_ack => ao_LL2_Out1_ack,
		In_rdy => ao_LL2_Out1_rdy,
		In_count => ao_LL2_Out1_count,
		-- Fanout Out
		Out_data => aof_LL2_Out1_data,
		Out_send => aof_LL2_Out1_send,
		Out_ack => aof_LL2_Out1_ack,
		Out_rdy => aof_LL2_Out1_rdy,
		Out_count => aof_LL2_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_LL1_iunzip_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_LL1_iunzip_Out1_data,
		In_send => ao_LL1_iunzip_Out1_send,
		In_ack => ao_LL1_iunzip_Out1_ack,
		In_rdy => ao_LL1_iunzip_Out1_rdy,
		In_count => ao_LL1_iunzip_Out1_count,
		-- Fanout Out
		Out_data => aof_LL1_iunzip_Out1_data,
		Out_send => aof_LL1_iunzip_Out1_send,
		Out_ack => aof_LL1_iunzip_Out1_ack,
		Out_rdy => aof_LL1_iunzip_Out1_rdy,
		Out_count => aof_LL1_iunzip_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	f_ao_LL1_iunzip_Out2 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_LL1_iunzip_Out2_data,
		In_send => ao_LL1_iunzip_Out2_send,
		In_ack => ao_LL1_iunzip_Out2_ack,
		In_rdy => ao_LL1_iunzip_Out2_rdy,
		In_count => ao_LL1_iunzip_Out2_count,
		-- Fanout Out
		Out_data => aof_LL1_iunzip_Out2_data,
		Out_send => aof_LL1_iunzip_Out2_send,
		Out_ack => aof_LL1_iunzip_Out2_ack,
		Out_rdy => aof_LL1_iunzip_Out2_rdy,
		Out_count => aof_LL1_iunzip_Out2_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_LL2_H_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_LL2_H_Out1_data,
		In_send => ao_LL2_H_Out1_send,
		In_ack => ao_LL2_H_Out1_ack,
		In_rdy => ao_LL2_H_Out1_rdy,
		In_count => ao_LL2_H_Out1_count,
		-- Fanout Out
		Out_data => aof_LL2_H_Out1_data,
		Out_send => aof_LL2_H_Out1_send,
		Out_ack => aof_LL2_H_Out1_ack,
		Out_rdy => aof_LL2_H_Out1_rdy,
		Out_count => aof_LL2_H_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_LL2_L_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_LL2_L_Out1_data,
		In_send => ao_LL2_L_Out1_send,
		In_ack => ao_LL2_L_Out1_ack,
		In_rdy => ao_LL2_L_Out1_rdy,
		In_count => ao_LL2_L_Out1_count,
		-- Fanout Out
		Out_data => aof_LL2_L_Out1_data,
		Out_send => aof_LL2_L_Out1_send,
		Out_ack => aof_LL2_L_Out1_ack,
		Out_rdy => aof_LL2_L_Out1_rdy,
		Out_count => aof_LL2_L_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_LL3_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_LL3_Out1_data,
		In_send => ao_LL3_Out1_send,
		In_ack => ao_LL3_Out1_ack,
		In_rdy => ao_LL3_Out1_rdy,
		In_count => ao_LL3_Out1_count,
		-- Fanout Out
		Out_data => aof_LL3_Out1_data,
		Out_send => aof_LL3_Out1_send,
		Out_ack => aof_LL3_Out1_ack,
		Out_rdy => aof_LL3_Out1_rdy,
		Out_count => aof_LL3_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_LL2_iunzip_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_LL2_iunzip_Out1_data,
		In_send => ao_LL2_iunzip_Out1_send,
		In_ack => ao_LL2_iunzip_Out1_ack,
		In_rdy => ao_LL2_iunzip_Out1_rdy,
		In_count => ao_LL2_iunzip_Out1_count,
		-- Fanout Out
		Out_data => aof_LL2_iunzip_Out1_data,
		Out_send => aof_LL2_iunzip_Out1_send,
		Out_ack => aof_LL2_iunzip_Out1_ack,
		Out_rdy => aof_LL2_iunzip_Out1_rdy,
		Out_count => aof_LL2_iunzip_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	f_ao_LL2_iunzip_Out2 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_LL2_iunzip_Out2_data,
		In_send => ao_LL2_iunzip_Out2_send,
		In_ack => ao_LL2_iunzip_Out2_ack,
		In_rdy => ao_LL2_iunzip_Out2_rdy,
		In_count => ao_LL2_iunzip_Out2_count,
		-- Fanout Out
		Out_data => aof_LL2_iunzip_Out2_data,
		Out_send => aof_LL2_iunzip_Out2_send,
		Out_ack => aof_LL2_iunzip_Out2_ack,
		Out_rdy => aof_LL2_iunzip_Out2_rdy,
		Out_count => aof_LL2_iunzip_Out2_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_LL3_H_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_LL3_H_Out1_data,
		In_send => ao_LL3_H_Out1_send,
		In_ack => ao_LL3_H_Out1_ack,
		In_rdy => ao_LL3_H_Out1_rdy,
		In_count => ao_LL3_H_Out1_count,
		-- Fanout Out
		Out_data => aof_LL3_H_Out1_data,
		Out_send => aof_LL3_H_Out1_send,
		Out_ack => aof_LL3_H_Out1_ack,
		Out_rdy => aof_LL3_H_Out1_rdy,
		Out_count => aof_LL3_H_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_LL3_L_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_LL3_L_Out1_data,
		In_send => ao_LL3_L_Out1_send,
		In_ack => ao_LL3_L_Out1_ack,
		In_rdy => ao_LL3_L_Out1_rdy,
		In_count => ao_LL3_L_Out1_count,
		-- Fanout Out
		Out_data => aof_LL3_L_Out1_data,
		Out_send => aof_LL3_L_Out1_send,
		Out_ack => aof_LL3_L_Out1_ack,
		Out_rdy => aof_LL3_L_Out1_rdy,
		Out_count => aof_LL3_L_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_image1_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_image1_Out1_data,
		In_send => ao_image1_Out1_send,
		In_ack => ao_image1_Out1_ack,
		In_rdy => ao_image1_Out1_rdy,
		In_count => ao_image1_Out1_count,
		-- Fanout Out
		Out_data => aof_image1_Out1_data,
		Out_send => aof_image1_Out1_send,
		Out_ack => aof_image1_Out1_ack,
		Out_rdy => aof_image1_Out1_rdy,
		Out_count => aof_image1_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_mapDia_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_mapDia_Out1_data,
		In_send => ao_mapDia_Out1_send,
		In_ack => ao_mapDia_Out1_ack,
		In_rdy => ao_mapDia_Out1_rdy,
		In_count => ao_mapDia_Out1_count,
		-- Fanout Out
		Out_data => aof_mapDia_Out1_data,
		Out_send => aof_mapDia_Out1_send,
		Out_ack => aof_mapDia_Out1_ack,
		Out_rdy => aof_mapDia_Out1_rdy,
		Out_count => aof_mapDia_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_mapFinal_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_mapFinal_Out1_data,
		In_send => ao_mapFinal_Out1_send,
		In_ack => ao_mapFinal_Out1_ack,
		In_rdy => ao_mapFinal_Out1_rdy,
		In_count => ao_mapFinal_Out1_count,
		-- Fanout Out
		Out_data => aof_mapFinal_Out1_data,
		Out_send => aof_mapFinal_Out1_send,
		Out_ack => aof_mapFinal_Out1_ack,
		Out_rdy => aof_mapFinal_Out1_rdy,
		Out_count => aof_mapFinal_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_mapVer_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_mapVer_Out1_data,
		In_send => ao_mapVer_Out1_send,
		In_ack => ao_mapVer_Out1_ack,
		In_rdy => ao_mapVer_Out1_rdy,
		In_count => ao_mapVer_Out1_count,
		-- Fanout Out
		Out_data => aof_mapVer_Out1_data,
		Out_send => aof_mapVer_Out1_send,
		Out_ack => aof_mapVer_Out1_ack,
		Out_rdy => aof_mapVer_Out1_rdy,
		Out_count => aof_mapVer_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_resized_HH1_xy_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_resized_HH1_xy_Out1_data,
		In_send => ao_resized_HH1_xy_Out1_send,
		In_ack => ao_resized_HH1_xy_Out1_ack,
		In_rdy => ao_resized_HH1_xy_Out1_rdy,
		In_count => ao_resized_HH1_xy_Out1_count,
		-- Fanout Out
		Out_data => aof_resized_HH1_xy_Out1_data,
		Out_send => aof_resized_HH1_xy_Out1_send,
		Out_ack => aof_resized_HH1_xy_Out1_ack,
		Out_rdy => aof_resized_HH1_xy_Out1_rdy,
		Out_count => aof_resized_HH1_xy_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_resized_HH1_xy_blurred_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_resized_HH1_xy_blurred_Out1_data,
		In_send => ao_resized_HH1_xy_blurred_Out1_send,
		In_ack => ao_resized_HH1_xy_blurred_Out1_ack,
		In_rdy => ao_resized_HH1_xy_blurred_Out1_rdy,
		In_count => ao_resized_HH1_xy_blurred_Out1_count,
		-- Fanout Out
		Out_data => aof_resized_HH1_xy_blurred_Out1_data,
		Out_send => aof_resized_HH1_xy_blurred_Out1_send,
		Out_ack => aof_resized_HH1_xy_blurred_Out1_ack,
		Out_rdy => aof_resized_HH1_xy_blurred_Out1_rdy,
		Out_count => aof_resized_HH1_xy_blurred_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_resized_HH2_xy_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_resized_HH2_xy_Out1_data,
		In_send => ao_resized_HH2_xy_Out1_send,
		In_ack => ao_resized_HH2_xy_Out1_ack,
		In_rdy => ao_resized_HH2_xy_Out1_rdy,
		In_count => ao_resized_HH2_xy_Out1_count,
		-- Fanout Out
		Out_data => aof_resized_HH2_xy_Out1_data,
		Out_send => aof_resized_HH2_xy_Out1_send,
		Out_ack => aof_resized_HH2_xy_Out1_ack,
		Out_rdy => aof_resized_HH2_xy_Out1_rdy,
		Out_count => aof_resized_HH2_xy_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_resized_HH2_xy_blurred_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_resized_HH2_xy_blurred_Out1_data,
		In_send => ao_resized_HH2_xy_blurred_Out1_send,
		In_ack => ao_resized_HH2_xy_blurred_Out1_ack,
		In_rdy => ao_resized_HH2_xy_blurred_Out1_rdy,
		In_count => ao_resized_HH2_xy_blurred_Out1_count,
		-- Fanout Out
		Out_data => aof_resized_HH2_xy_blurred_Out1_data,
		Out_send => aof_resized_HH2_xy_blurred_Out1_send,
		Out_ack => aof_resized_HH2_xy_blurred_Out1_ack,
		Out_rdy => aof_resized_HH2_xy_blurred_Out1_rdy,
		Out_count => aof_resized_HH2_xy_blurred_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_resized_HH3_xy_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_resized_HH3_xy_Out1_data,
		In_send => ao_resized_HH3_xy_Out1_send,
		In_ack => ao_resized_HH3_xy_Out1_ack,
		In_rdy => ao_resized_HH3_xy_Out1_rdy,
		In_count => ao_resized_HH3_xy_Out1_count,
		-- Fanout Out
		Out_data => aof_resized_HH3_xy_Out1_data,
		Out_send => aof_resized_HH3_xy_Out1_send,
		Out_ack => aof_resized_HH3_xy_Out1_ack,
		Out_rdy => aof_resized_HH3_xy_Out1_rdy,
		Out_count => aof_resized_HH3_xy_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_resized_HH3_xy_blurred_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_resized_HH3_xy_blurred_Out1_data,
		In_send => ao_resized_HH3_xy_blurred_Out1_send,
		In_ack => ao_resized_HH3_xy_blurred_Out1_ack,
		In_rdy => ao_resized_HH3_xy_blurred_Out1_rdy,
		In_count => ao_resized_HH3_xy_blurred_Out1_count,
		-- Fanout Out
		Out_data => aof_resized_HH3_xy_blurred_Out1_data,
		Out_send => aof_resized_HH3_xy_blurred_Out1_send,
		Out_ack => aof_resized_HH3_xy_blurred_Out1_ack,
		Out_rdy => aof_resized_HH3_xy_blurred_Out1_rdy,
		Out_count => aof_resized_HH3_xy_blurred_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_resized_LH1_xy_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_resized_LH1_xy_Out1_data,
		In_send => ao_resized_LH1_xy_Out1_send,
		In_ack => ao_resized_LH1_xy_Out1_ack,
		In_rdy => ao_resized_LH1_xy_Out1_rdy,
		In_count => ao_resized_LH1_xy_Out1_count,
		-- Fanout Out
		Out_data => aof_resized_LH1_xy_Out1_data,
		Out_send => aof_resized_LH1_xy_Out1_send,
		Out_ack => aof_resized_LH1_xy_Out1_ack,
		Out_rdy => aof_resized_LH1_xy_Out1_rdy,
		Out_count => aof_resized_LH1_xy_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_resized_LH1_xy_blurred_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_resized_LH1_xy_blurred_Out1_data,
		In_send => ao_resized_LH1_xy_blurred_Out1_send,
		In_ack => ao_resized_LH1_xy_blurred_Out1_ack,
		In_rdy => ao_resized_LH1_xy_blurred_Out1_rdy,
		In_count => ao_resized_LH1_xy_blurred_Out1_count,
		-- Fanout Out
		Out_data => aof_resized_LH1_xy_blurred_Out1_data,
		Out_send => aof_resized_LH1_xy_blurred_Out1_send,
		Out_ack => aof_resized_LH1_xy_blurred_Out1_ack,
		Out_rdy => aof_resized_LH1_xy_blurred_Out1_rdy,
		Out_count => aof_resized_LH1_xy_blurred_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_resized_LH2_xy_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_resized_LH2_xy_Out1_data,
		In_send => ao_resized_LH2_xy_Out1_send,
		In_ack => ao_resized_LH2_xy_Out1_ack,
		In_rdy => ao_resized_LH2_xy_Out1_rdy,
		In_count => ao_resized_LH2_xy_Out1_count,
		-- Fanout Out
		Out_data => aof_resized_LH2_xy_Out1_data,
		Out_send => aof_resized_LH2_xy_Out1_send,
		Out_ack => aof_resized_LH2_xy_Out1_ack,
		Out_rdy => aof_resized_LH2_xy_Out1_rdy,
		Out_count => aof_resized_LH2_xy_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_resized_LH2_xy_blurred_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_resized_LH2_xy_blurred_Out1_data,
		In_send => ao_resized_LH2_xy_blurred_Out1_send,
		In_ack => ao_resized_LH2_xy_blurred_Out1_ack,
		In_rdy => ao_resized_LH2_xy_blurred_Out1_rdy,
		In_count => ao_resized_LH2_xy_blurred_Out1_count,
		-- Fanout Out
		Out_data => aof_resized_LH2_xy_blurred_Out1_data,
		Out_send => aof_resized_LH2_xy_blurred_Out1_send,
		Out_ack => aof_resized_LH2_xy_blurred_Out1_ack,
		Out_rdy => aof_resized_LH2_xy_blurred_Out1_rdy,
		Out_count => aof_resized_LH2_xy_blurred_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_resized_LH3_xy_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_resized_LH3_xy_Out1_data,
		In_send => ao_resized_LH3_xy_Out1_send,
		In_ack => ao_resized_LH3_xy_Out1_ack,
		In_rdy => ao_resized_LH3_xy_Out1_rdy,
		In_count => ao_resized_LH3_xy_Out1_count,
		-- Fanout Out
		Out_data => aof_resized_LH3_xy_Out1_data,
		Out_send => aof_resized_LH3_xy_Out1_send,
		Out_ack => aof_resized_LH3_xy_Out1_ack,
		Out_rdy => aof_resized_LH3_xy_Out1_rdy,
		Out_count => aof_resized_LH3_xy_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));
	
	f_ao_resized_LH3_xy_blurred_Out1 : entity SystemBuilder.Fanout(behavioral)
	generic map (fanout => 1, width => 16)
	port map(
		-- Fanout In
		In_data => ao_resized_LH3_xy_blurred_Out1_data,
		In_send => ao_resized_LH3_xy_blurred_Out1_send,
		In_ack => ao_resized_LH3_xy_blurred_Out1_ack,
		In_rdy => ao_resized_LH3_xy_blurred_Out1_rdy,
		In_count => ao_resized_LH3_xy_blurred_Out1_count,
		-- Fanout Out
		Out_data => aof_resized_LH3_xy_blurred_Out1_data,
		Out_send => aof_resized_LH3_xy_blurred_Out1_send,
		Out_ack => aof_resized_LH3_xy_blurred_Out1_ack,
		Out_rdy => aof_resized_LH3_xy_blurred_Out1_rdy,
		Out_count => aof_resized_LH3_xy_blurred_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0));

	-- --------------------------------------------------------------------------
	-- Queues
	-- --------------------------------------------------------------------------
	q_ai_HH1_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_HH1_In1_data,
		Out_send => ai_HH1_In1_send,
		Out_ack => ai_HH1_In1_ack,
		Out_count => ai_HH1_In1_count,
		-- Queue In
		In_data => aof_LL1_H_iunzipFilter2D_Out2_data,
		In_send => aof_LL1_H_iunzipFilter2D_Out2_send(0),
		In_ack => aof_LL1_H_iunzipFilter2D_Out2_ack(0),
		In_rdy => aof_LL1_H_iunzipFilter2D_Out2_rdy(0),
		In_count => aof_LL1_H_iunzipFilter2D_Out2_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_LL1_H_iunzipFilter2D_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_LL1_H_iunzipFilter2D_In1_data,
		Out_send => ai_LL1_H_iunzipFilter2D_In1_send,
		Out_ack => ai_LL1_H_iunzipFilter2D_In1_ack,
		Out_count => ai_LL1_H_iunzipFilter2D_In1_count,
		-- Queue In
		In_data => aof_LL1_H_Out1_data,
		In_send => aof_LL1_H_Out1_send(0),
		In_ack => aof_LL1_H_Out1_ack(0),
		In_rdy => aof_LL1_H_Out1_rdy(0),
		In_count => aof_LL1_H_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_HH2_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_HH2_In1_data,
		Out_send => ai_HH2_In1_send,
		Out_ack => ai_HH2_In1_ack,
		Out_count => ai_HH2_In1_count,
		-- Queue In
		In_data => aof_LL2_H_iunzipFilter2D_Out2_data,
		In_send => aof_LL2_H_iunzipFilter2D_Out2_send(0),
		In_ack => aof_LL2_H_iunzipFilter2D_Out2_ack(0),
		In_rdy => aof_LL2_H_iunzipFilter2D_Out2_rdy(0),
		In_count => aof_LL2_H_iunzipFilter2D_Out2_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_LL2_H_iunzipFilter2D_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_LL2_H_iunzipFilter2D_In1_data,
		Out_send => ai_LL2_H_iunzipFilter2D_In1_send,
		Out_ack => ai_LL2_H_iunzipFilter2D_In1_ack,
		Out_count => ai_LL2_H_iunzipFilter2D_In1_count,
		-- Queue In
		In_data => aof_LL2_H_Out1_data,
		In_send => aof_LL2_H_Out1_send(0),
		In_ack => aof_LL2_H_Out1_ack(0),
		In_rdy => aof_LL2_H_Out1_rdy(0),
		In_count => aof_LL2_H_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_HH3_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_HH3_In1_data,
		Out_send => ai_HH3_In1_send,
		Out_ack => ai_HH3_In1_ack,
		Out_count => ai_HH3_In1_count,
		-- Queue In
		In_data => aof_LL3_H_iunzipFilter2D_Out2_data,
		In_send => aof_LL3_H_iunzipFilter2D_Out2_send(0),
		In_ack => aof_LL3_H_iunzipFilter2D_Out2_ack(0),
		In_rdy => aof_LL3_H_iunzipFilter2D_Out2_rdy(0),
		In_count => aof_LL3_H_iunzipFilter2D_Out2_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_LL3_H_iunzipFilter2D_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_LL3_H_iunzipFilter2D_In1_data,
		Out_send => ai_LL3_H_iunzipFilter2D_In1_send,
		Out_ack => ai_LL3_H_iunzipFilter2D_In1_ack,
		Out_count => ai_LL3_H_iunzipFilter2D_In1_count,
		-- Queue In
		In_data => aof_LL3_H_Out1_data,
		In_send => aof_LL3_H_Out1_send(0),
		In_ack => aof_LL3_H_Out1_ack(0),
		In_rdy => aof_LL3_H_Out1_rdy(0),
		In_count => aof_LL3_H_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_HL1_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_HL1_In1_data,
		Out_send => ai_HL1_In1_send,
		Out_ack => ai_HL1_In1_ack,
		Out_count => ai_HL1_In1_count,
		-- Queue In
		In_data => aof_LL1_H_iunzipFilter2D_Out1_data,
		In_send => aof_LL1_H_iunzipFilter2D_Out1_send(0),
		In_ack => aof_LL1_H_iunzipFilter2D_Out1_ack(0),
		In_rdy => aof_LL1_H_iunzipFilter2D_Out1_rdy(0),
		In_count => aof_LL1_H_iunzipFilter2D_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_HL2_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_HL2_In1_data,
		Out_send => ai_HL2_In1_send,
		Out_ack => ai_HL2_In1_ack,
		Out_count => ai_HL2_In1_count,
		-- Queue In
		In_data => aof_LL2_H_iunzipFilter2D_Out1_data,
		In_send => aof_LL2_H_iunzipFilter2D_Out1_send(0),
		In_ack => aof_LL2_H_iunzipFilter2D_Out1_ack(0),
		In_rdy => aof_LL2_H_iunzipFilter2D_Out1_rdy(0),
		In_count => aof_LL2_H_iunzipFilter2D_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_HL3_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_HL3_In1_data,
		Out_send => ai_HL3_In1_send,
		Out_ack => ai_HL3_In1_ack,
		Out_count => ai_HL3_In1_count,
		-- Queue In
		In_data => aof_LL3_H_iunzipFilter2D_Out1_data,
		In_send => aof_LL3_H_iunzipFilter2D_Out1_send(0),
		In_ack => aof_LL3_H_iunzipFilter2D_Out1_ack(0),
		In_rdy => aof_LL3_H_iunzipFilter2D_Out1_rdy(0),
		In_count => aof_LL3_H_iunzipFilter2D_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_LH1_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_LH1_In1_data,
		Out_send => ai_LH1_In1_send,
		Out_ack => ai_LH1_In1_ack,
		Out_count => ai_LH1_In1_count,
		-- Queue In
		In_data => aof_LL1_L_iunzipFilter2D_Out2_data,
		In_send => aof_LL1_L_iunzipFilter2D_Out2_send(0),
		In_ack => aof_LL1_L_iunzipFilter2D_Out2_ack(0),
		In_rdy => aof_LL1_L_iunzipFilter2D_Out2_rdy(0),
		In_count => aof_LL1_L_iunzipFilter2D_Out2_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_LL1_L_iunzipFilter2D_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_LL1_L_iunzipFilter2D_In1_data,
		Out_send => ai_LL1_L_iunzipFilter2D_In1_send,
		Out_ack => ai_LL1_L_iunzipFilter2D_In1_ack,
		Out_count => ai_LL1_L_iunzipFilter2D_In1_count,
		-- Queue In
		In_data => aof_LL1_L_Out1_data,
		In_send => aof_LL1_L_Out1_send(0),
		In_ack => aof_LL1_L_Out1_ack(0),
		In_rdy => aof_LL1_L_Out1_rdy(0),
		In_count => aof_LL1_L_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_LH2_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_LH2_In1_data,
		Out_send => ai_LH2_In1_send,
		Out_ack => ai_LH2_In1_ack,
		Out_count => ai_LH2_In1_count,
		-- Queue In
		In_data => aof_LL2_L_iunzipFilter2D_Out2_data,
		In_send => aof_LL2_L_iunzipFilter2D_Out2_send(0),
		In_ack => aof_LL2_L_iunzipFilter2D_Out2_ack(0),
		In_rdy => aof_LL2_L_iunzipFilter2D_Out2_rdy(0),
		In_count => aof_LL2_L_iunzipFilter2D_Out2_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_LL2_L_iunzipFilter2D_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_LL2_L_iunzipFilter2D_In1_data,
		Out_send => ai_LL2_L_iunzipFilter2D_In1_send,
		Out_ack => ai_LL2_L_iunzipFilter2D_In1_ack,
		Out_count => ai_LL2_L_iunzipFilter2D_In1_count,
		-- Queue In
		In_data => aof_LL2_L_Out1_data,
		In_send => aof_LL2_L_Out1_send(0),
		In_ack => aof_LL2_L_Out1_ack(0),
		In_rdy => aof_LL2_L_Out1_rdy(0),
		In_count => aof_LL2_L_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_LH3_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_LH3_In1_data,
		Out_send => ai_LH3_In1_send,
		Out_ack => ai_LH3_In1_ack,
		Out_count => ai_LH3_In1_count,
		-- Queue In
		In_data => aof_LL3_L_iunzipFilter2D_Out2_data,
		In_send => aof_LL3_L_iunzipFilter2D_Out2_send(0),
		In_ack => aof_LL3_L_iunzipFilter2D_Out2_ack(0),
		In_rdy => aof_LL3_L_iunzipFilter2D_Out2_rdy(0),
		In_count => aof_LL3_L_iunzipFilter2D_Out2_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_LL3_L_iunzipFilter2D_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_LL3_L_iunzipFilter2D_In1_data,
		Out_send => ai_LL3_L_iunzipFilter2D_In1_send,
		Out_ack => ai_LL3_L_iunzipFilter2D_In1_ack,
		Out_count => ai_LL3_L_iunzipFilter2D_In1_count,
		-- Queue In
		In_data => aof_LL3_L_Out1_data,
		In_send => aof_LL3_L_Out1_send(0),
		In_ack => aof_LL3_L_Out1_ack(0),
		In_rdy => aof_LL3_L_Out1_rdy(0),
		In_count => aof_LL3_L_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_LL1_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_LL1_In1_data,
		Out_send => ai_LL1_In1_send,
		Out_ack => ai_LL1_In1_ack,
		Out_count => ai_LL1_In1_count,
		-- Queue In
		In_data => aof_LL1_L_iunzipFilter2D_Out1_data,
		In_send => aof_LL1_L_iunzipFilter2D_Out1_send(0),
		In_ack => aof_LL1_L_iunzipFilter2D_Out1_ack(0),
		In_rdy => aof_LL1_L_iunzipFilter2D_Out1_rdy(0),
		In_count => aof_LL1_L_iunzipFilter2D_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_LL1_H_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_LL1_H_In1_data,
		Out_send => ai_LL1_H_In1_send,
		Out_ack => ai_LL1_H_In1_ack,
		Out_count => ai_LL1_H_In1_count,
		-- Queue In
		In_data => aof_image1_iunzip_Out2_data,
		In_send => aof_image1_iunzip_Out2_send(0),
		In_ack => aof_image1_iunzip_Out2_ack(0),
		In_rdy => aof_image1_iunzip_Out2_rdy(0),
		In_count => aof_image1_iunzip_Out2_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_image1_iunzip_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_image1_iunzip_In1_data,
		Out_send => ai_image1_iunzip_In1_send,
		Out_ack => ai_image1_iunzip_In1_ack,
		Out_count => ai_image1_iunzip_In1_count,
		-- Queue In
		In_data => aof_image1_Out1_data,
		In_send => aof_image1_Out1_send(0),
		In_ack => aof_image1_Out1_ack(0),
		In_rdy => aof_image1_Out1_rdy(0),
		In_count => aof_image1_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_LL1_L_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_LL1_L_In1_data,
		Out_send => ai_LL1_L_In1_send,
		Out_ack => ai_LL1_L_In1_ack,
		Out_count => ai_LL1_L_In1_count,
		-- Queue In
		In_data => aof_image1_iunzip_Out1_data,
		In_send => aof_image1_iunzip_Out1_send(0),
		In_ack => aof_image1_iunzip_Out1_ack(0),
		In_rdy => aof_image1_iunzip_Out1_rdy(0),
		In_count => aof_image1_iunzip_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_LL2_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_LL2_In1_data,
		Out_send => ai_LL2_In1_send,
		Out_ack => ai_LL2_In1_ack,
		Out_count => ai_LL2_In1_count,
		-- Queue In
		In_data => aof_LL2_L_iunzipFilter2D_Out1_data,
		In_send => aof_LL2_L_iunzipFilter2D_Out1_send(0),
		In_ack => aof_LL2_L_iunzipFilter2D_Out1_ack(0),
		In_rdy => aof_LL2_L_iunzipFilter2D_Out1_rdy(0),
		In_count => aof_LL2_L_iunzipFilter2D_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_LL2_H_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_LL2_H_In1_data,
		Out_send => ai_LL2_H_In1_send,
		Out_ack => ai_LL2_H_In1_ack,
		Out_count => ai_LL2_H_In1_count,
		-- Queue In
		In_data => aof_LL1_iunzip_Out2_data,
		In_send => aof_LL1_iunzip_Out2_send(0),
		In_ack => aof_LL1_iunzip_Out2_ack(0),
		In_rdy => aof_LL1_iunzip_Out2_rdy(0),
		In_count => aof_LL1_iunzip_Out2_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_LL1_iunzip_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_LL1_iunzip_In1_data,
		Out_send => ai_LL1_iunzip_In1_send,
		Out_ack => ai_LL1_iunzip_In1_ack,
		Out_count => ai_LL1_iunzip_In1_count,
		-- Queue In
		In_data => aof_LL1_Out1_data,
		In_send => aof_LL1_Out1_send(0),
		In_ack => aof_LL1_Out1_ack(0),
		In_rdy => aof_LL1_Out1_rdy(0),
		In_count => aof_LL1_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_LL2_L_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_LL2_L_In1_data,
		Out_send => ai_LL2_L_In1_send,
		Out_ack => ai_LL2_L_In1_ack,
		Out_count => ai_LL2_L_In1_count,
		-- Queue In
		In_data => aof_LL1_iunzip_Out1_data,
		In_send => aof_LL1_iunzip_Out1_send(0),
		In_ack => aof_LL1_iunzip_Out1_ack(0),
		In_rdy => aof_LL1_iunzip_Out1_rdy(0),
		In_count => aof_LL1_iunzip_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_LL3_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_LL3_In1_data,
		Out_send => ai_LL3_In1_send,
		Out_ack => ai_LL3_In1_ack,
		Out_count => ai_LL3_In1_count,
		-- Queue In
		In_data => aof_LL3_L_iunzipFilter2D_Out1_data,
		In_send => aof_LL3_L_iunzipFilter2D_Out1_send(0),
		In_ack => aof_LL3_L_iunzipFilter2D_Out1_ack(0),
		In_rdy => aof_LL3_L_iunzipFilter2D_Out1_rdy(0),
		In_count => aof_LL3_L_iunzipFilter2D_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_LL3_H_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_LL3_H_In1_data,
		Out_send => ai_LL3_H_In1_send,
		Out_ack => ai_LL3_H_In1_ack,
		Out_count => ai_LL3_H_In1_count,
		-- Queue In
		In_data => aof_LL2_iunzip_Out2_data,
		In_send => aof_LL2_iunzip_Out2_send(0),
		In_ack => aof_LL2_iunzip_Out2_ack(0),
		In_rdy => aof_LL2_iunzip_Out2_rdy(0),
		In_count => aof_LL2_iunzip_Out2_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_LL2_iunzip_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_LL2_iunzip_In1_data,
		Out_send => ai_LL2_iunzip_In1_send,
		Out_ack => ai_LL2_iunzip_In1_ack,
		Out_count => ai_LL2_iunzip_In1_count,
		-- Queue In
		In_data => aof_LL2_Out1_data,
		In_send => aof_LL2_Out1_send(0),
		In_ack => aof_LL2_Out1_ack(0),
		In_rdy => aof_LL2_Out1_rdy(0),
		In_count => aof_LL2_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_LL3_L_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_LL3_L_In1_data,
		Out_send => ai_LL3_L_In1_send,
		Out_ack => ai_LL3_L_In1_ack,
		Out_count => ai_LL3_L_In1_count,
		-- Queue In
		In_data => aof_LL2_iunzip_Out1_data,
		In_send => aof_LL2_iunzip_Out1_send(0),
		In_ack => aof_LL2_iunzip_Out1_ack(0),
		In_rdy => aof_LL2_iunzip_Out1_rdy(0),
		In_count => aof_LL2_iunzip_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_image1_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_image1_In1_data,
		Out_send => ai_image1_In1_send,
		Out_ack => ai_image1_In1_ack,
		Out_count => ai_image1_In1_count,
		-- Queue In
		In_data => nif_In_data,
		In_send => nif_In_send(0),
		In_ack => nif_In_ack(0),
		In_rdy => nif_In_rdy(0),
		In_count => nif_In_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_mapDia_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_mapDia_In1_data,
		Out_send => ai_mapDia_In1_send,
		Out_ack => ai_mapDia_In1_ack,
		Out_count => ai_mapDia_In1_count,
		-- Queue In
		In_data => aof_resized_HH1_xy_Out1_data,
		In_send => aof_resized_HH1_xy_Out1_send(0),
		In_ack => aof_resized_HH1_xy_Out1_ack(0),
		In_rdy => aof_resized_HH1_xy_Out1_rdy(0),
		In_count => aof_resized_HH1_xy_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_mapDia_In2 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_mapDia_In2_data,
		Out_send => ai_mapDia_In2_send,
		Out_ack => ai_mapDia_In2_ack,
		Out_count => ai_mapDia_In2_count,
		-- Queue In
		In_data => aof_resized_HH2_xy_Out1_data,
		In_send => aof_resized_HH2_xy_Out1_send(0),
		In_ack => aof_resized_HH2_xy_Out1_ack(0),
		In_rdy => aof_resized_HH2_xy_Out1_rdy(0),
		In_count => aof_resized_HH2_xy_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_mapDia_In3 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_mapDia_In3_data,
		Out_send => ai_mapDia_In3_send,
		Out_ack => ai_mapDia_In3_ack,
		Out_count => ai_mapDia_In3_count,
		-- Queue In
		In_data => aof_resized_HH3_xy_Out1_data,
		In_send => aof_resized_HH3_xy_Out1_send(0),
		In_ack => aof_resized_HH3_xy_Out1_ack(0),
		In_rdy => aof_resized_HH3_xy_Out1_rdy(0),
		In_count => aof_resized_HH3_xy_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_mapFinal_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_mapFinal_In1_data,
		Out_send => ai_mapFinal_In1_send,
		Out_ack => ai_mapFinal_In1_ack,
		Out_count => ai_mapFinal_In1_count,
		-- Queue In
		In_data => aof_mapVer_Out1_data,
		In_send => aof_mapVer_Out1_send(0),
		In_ack => aof_mapVer_Out1_ack(0),
		In_rdy => aof_mapVer_Out1_rdy(0),
		In_count => aof_mapVer_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_mapFinal_In2 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_mapFinal_In2_data,
		Out_send => ai_mapFinal_In2_send,
		Out_ack => ai_mapFinal_In2_ack,
		Out_count => ai_mapFinal_In2_count,
		-- Queue In
		In_data => aof_mapDia_Out1_data,
		In_send => aof_mapDia_Out1_send(0),
		In_ack => aof_mapDia_Out1_ack(0),
		In_rdy => aof_mapDia_Out1_rdy(0),
		In_count => aof_mapDia_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_mapVer_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_mapVer_In1_data,
		Out_send => ai_mapVer_In1_send,
		Out_ack => ai_mapVer_In1_ack,
		Out_count => ai_mapVer_In1_count,
		-- Queue In
		In_data => aof_resized_LH1_xy_Out1_data,
		In_send => aof_resized_LH1_xy_Out1_send(0),
		In_ack => aof_resized_LH1_xy_Out1_ack(0),
		In_rdy => aof_resized_LH1_xy_Out1_rdy(0),
		In_count => aof_resized_LH1_xy_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_mapVer_In2 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_mapVer_In2_data,
		Out_send => ai_mapVer_In2_send,
		Out_ack => ai_mapVer_In2_ack,
		Out_count => ai_mapVer_In2_count,
		-- Queue In
		In_data => aof_resized_LH2_xy_Out1_data,
		In_send => aof_resized_LH2_xy_Out1_send(0),
		In_ack => aof_resized_LH2_xy_Out1_ack(0),
		In_rdy => aof_resized_LH2_xy_Out1_rdy(0),
		In_count => aof_resized_LH2_xy_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_mapVer_In3 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_mapVer_In3_data,
		Out_send => ai_mapVer_In3_send,
		Out_ack => ai_mapVer_In3_ack,
		Out_count => ai_mapVer_In3_count,
		-- Queue In
		In_data => aof_resized_LH3_xy_Out1_data,
		In_send => aof_resized_LH3_xy_Out1_send(0),
		In_ack => aof_resized_LH3_xy_Out1_ack(0),
		In_rdy => aof_resized_LH3_xy_Out1_rdy(0),
		In_count => aof_resized_LH3_xy_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_no_Out : entity SystemBuilder.Queue(behavioral)
	generic map (length => 64, width => 16)
	port map(
		-- Queue Out
		Out_data => no_Out_data,
		Out_send => no_Out_send,
		Out_ack => no_Out_ack,
		Out_count => no_Out_count,
		-- Queue In
		In_data => aof_mapFinal_Out1_data,
		In_send => aof_mapFinal_Out1_send(0),
		In_ack => aof_mapFinal_Out1_ack(0),
		In_rdy => aof_mapFinal_Out1_rdy(0),
		In_count => aof_mapFinal_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_resized_HH1_xy_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_resized_HH1_xy_In1_data,
		Out_send => ai_resized_HH1_xy_In1_send,
		Out_ack => ai_resized_HH1_xy_In1_ack,
		Out_count => ai_resized_HH1_xy_In1_count,
		-- Queue In
		In_data => aof_resized_HH1_xy_blurred_Out1_data,
		In_send => aof_resized_HH1_xy_blurred_Out1_send(0),
		In_ack => aof_resized_HH1_xy_blurred_Out1_ack(0),
		In_rdy => aof_resized_HH1_xy_blurred_Out1_rdy(0),
		In_count => aof_resized_HH1_xy_blurred_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_resized_HH1_xy_blurred_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_resized_HH1_xy_blurred_In1_data,
		Out_send => ai_resized_HH1_xy_blurred_In1_send,
		Out_ack => ai_resized_HH1_xy_blurred_In1_ack,
		Out_count => ai_resized_HH1_xy_blurred_In1_count,
		-- Queue In
		In_data => aof_HH1_Out1_data,
		In_send => aof_HH1_Out1_send(0),
		In_ack => aof_HH1_Out1_ack(0),
		In_rdy => aof_HH1_Out1_rdy(0),
		In_count => aof_HH1_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_resized_HH2_xy_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_resized_HH2_xy_In1_data,
		Out_send => ai_resized_HH2_xy_In1_send,
		Out_ack => ai_resized_HH2_xy_In1_ack,
		Out_count => ai_resized_HH2_xy_In1_count,
		-- Queue In
		In_data => aof_resized_HH2_xy_blurred_Out1_data,
		In_send => aof_resized_HH2_xy_blurred_Out1_send(0),
		In_ack => aof_resized_HH2_xy_blurred_Out1_ack(0),
		In_rdy => aof_resized_HH2_xy_blurred_Out1_rdy(0),
		In_count => aof_resized_HH2_xy_blurred_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_resized_HH2_xy_blurred_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_resized_HH2_xy_blurred_In1_data,
		Out_send => ai_resized_HH2_xy_blurred_In1_send,
		Out_ack => ai_resized_HH2_xy_blurred_In1_ack,
		Out_count => ai_resized_HH2_xy_blurred_In1_count,
		-- Queue In
		In_data => aof_HH2_Out1_data,
		In_send => aof_HH2_Out1_send(0),
		In_ack => aof_HH2_Out1_ack(0),
		In_rdy => aof_HH2_Out1_rdy(0),
		In_count => aof_HH2_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_resized_HH3_xy_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_resized_HH3_xy_In1_data,
		Out_send => ai_resized_HH3_xy_In1_send,
		Out_ack => ai_resized_HH3_xy_In1_ack,
		Out_count => ai_resized_HH3_xy_In1_count,
		-- Queue In
		In_data => aof_resized_HH3_xy_blurred_Out1_data,
		In_send => aof_resized_HH3_xy_blurred_Out1_send(0),
		In_ack => aof_resized_HH3_xy_blurred_Out1_ack(0),
		In_rdy => aof_resized_HH3_xy_blurred_Out1_rdy(0),
		In_count => aof_resized_HH3_xy_blurred_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_resized_HH3_xy_blurred_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_resized_HH3_xy_blurred_In1_data,
		Out_send => ai_resized_HH3_xy_blurred_In1_send,
		Out_ack => ai_resized_HH3_xy_blurred_In1_ack,
		Out_count => ai_resized_HH3_xy_blurred_In1_count,
		-- Queue In
		In_data => aof_HH3_Out1_data,
		In_send => aof_HH3_Out1_send(0),
		In_ack => aof_HH3_Out1_ack(0),
		In_rdy => aof_HH3_Out1_rdy(0),
		In_count => aof_HH3_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_resized_LH1_xy_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_resized_LH1_xy_In1_data,
		Out_send => ai_resized_LH1_xy_In1_send,
		Out_ack => ai_resized_LH1_xy_In1_ack,
		Out_count => ai_resized_LH1_xy_In1_count,
		-- Queue In
		In_data => aof_resized_LH1_xy_blurred_Out1_data,
		In_send => aof_resized_LH1_xy_blurred_Out1_send(0),
		In_ack => aof_resized_LH1_xy_blurred_Out1_ack(0),
		In_rdy => aof_resized_LH1_xy_blurred_Out1_rdy(0),
		In_count => aof_resized_LH1_xy_blurred_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_resized_LH1_xy_blurred_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_resized_LH1_xy_blurred_In1_data,
		Out_send => ai_resized_LH1_xy_blurred_In1_send,
		Out_ack => ai_resized_LH1_xy_blurred_In1_ack,
		Out_count => ai_resized_LH1_xy_blurred_In1_count,
		-- Queue In
		In_data => aof_LH1_Out1_data,
		In_send => aof_LH1_Out1_send(0),
		In_ack => aof_LH1_Out1_ack(0),
		In_rdy => aof_LH1_Out1_rdy(0),
		In_count => aof_LH1_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_resized_LH2_xy_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_resized_LH2_xy_In1_data,
		Out_send => ai_resized_LH2_xy_In1_send,
		Out_ack => ai_resized_LH2_xy_In1_ack,
		Out_count => ai_resized_LH2_xy_In1_count,
		-- Queue In
		In_data => aof_resized_LH2_xy_blurred_Out1_data,
		In_send => aof_resized_LH2_xy_blurred_Out1_send(0),
		In_ack => aof_resized_LH2_xy_blurred_Out1_ack(0),
		In_rdy => aof_resized_LH2_xy_blurred_Out1_rdy(0),
		In_count => aof_resized_LH2_xy_blurred_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_resized_LH2_xy_blurred_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_resized_LH2_xy_blurred_In1_data,
		Out_send => ai_resized_LH2_xy_blurred_In1_send,
		Out_ack => ai_resized_LH2_xy_blurred_In1_ack,
		Out_count => ai_resized_LH2_xy_blurred_In1_count,
		-- Queue In
		In_data => aof_LH2_Out1_data,
		In_send => aof_LH2_Out1_send(0),
		In_ack => aof_LH2_Out1_ack(0),
		In_rdy => aof_LH2_Out1_rdy(0),
		In_count => aof_LH2_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_resized_LH3_xy_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_resized_LH3_xy_In1_data,
		Out_send => ai_resized_LH3_xy_In1_send,
		Out_ack => ai_resized_LH3_xy_In1_ack,
		Out_count => ai_resized_LH3_xy_In1_count,
		-- Queue In
		In_data => aof_resized_LH3_xy_blurred_Out1_data,
		In_send => aof_resized_LH3_xy_blurred_Out1_send(0),
		In_ack => aof_resized_LH3_xy_blurred_Out1_ack(0),
		In_rdy => aof_resized_LH3_xy_blurred_Out1_rdy(0),
		In_count => aof_resized_LH3_xy_blurred_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_ai_resized_LH3_xy_blurred_In1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 4, width => 16)
	port map(
		-- Queue Out
		Out_data => ai_resized_LH3_xy_blurred_In1_data,
		Out_send => ai_resized_LH3_xy_blurred_In1_send,
		Out_ack => ai_resized_LH3_xy_blurred_In1_ack,
		Out_count => ai_resized_LH3_xy_blurred_In1_count,
		-- Queue In
		In_data => aof_LH3_Out1_data,
		In_send => aof_LH3_Out1_send(0),
		In_ack => aof_LH3_Out1_ack(0),
		In_rdy => aof_LH3_Out1_rdy(0),
		In_count => aof_LH3_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_no_dummy1 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 64, width => 16)
	port map(
		-- Queue Out
		Out_data => no_dummy1_data,
		Out_send => no_dummy1_send,
		Out_ack => no_dummy1_ack,
		Out_count => no_dummy1_count,
		-- Queue In
		In_data => aof_HL1_Out1_data,
		In_send => aof_HL1_Out1_send(0),
		In_ack => aof_HL1_Out1_ack(0),
		In_rdy => aof_HL1_Out1_rdy(0),
		In_count => aof_HL1_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_no_dummy2 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 64, width => 16)
	port map(
		-- Queue Out
		Out_data => no_dummy2_data,
		Out_send => no_dummy2_send,
		Out_ack => no_dummy2_ack,
		Out_count => no_dummy2_count,
		-- Queue In
		In_data => aof_HL2_Out1_data,
		In_send => aof_HL2_Out1_send(0),
		In_ack => aof_HL2_Out1_ack(0),
		In_rdy => aof_HL2_Out1_rdy(0),
		In_count => aof_HL2_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_no_dummy3 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 64, width => 16)
	port map(
		-- Queue Out
		Out_data => no_dummy3_data,
		Out_send => no_dummy3_send,
		Out_ack => no_dummy3_ack,
		Out_count => no_dummy3_count,
		-- Queue In
		In_data => aof_HL3_Out1_data,
		In_send => aof_HL3_Out1_send(0),
		In_ack => aof_HL3_Out1_ack(0),
		In_rdy => aof_HL3_Out1_rdy(0),
		In_count => aof_HL3_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);
	
	q_no_dummy4 : entity SystemBuilder.Queue(behavioral)
	generic map (length => 64, width => 16)
	port map(
		-- Queue Out
		Out_data => no_dummy4_data,
		Out_send => no_dummy4_send,
		Out_ack => no_dummy4_ack,
		Out_count => no_dummy4_count,
		-- Queue In
		In_data => aof_LL3_Out1_data,
		In_send => aof_LL3_Out1_send(0),
		In_ack => aof_LL3_Out1_ack(0),
		In_rdy => aof_LL3_Out1_rdy(0),
		In_count => aof_LL3_Out1_count,
		-- Clock & Reset
		clk => clocks(0),
		reset => resets(0)
	);

	-- --------------------------------------------------------------------------
	-- Network port(s) instantiation
	-- --------------------------------------------------------------------------
	
	-- Output Port(s) Instantiation
	Out_data <= no_Out_data;
	Out_send <= no_Out_send;
	no_Out_ack <= Out_ack;
	no_Out_rdy <= Out_rdy;
	Out_count <= no_Out_count;
	dummy1_data <= no_dummy1_data;
	dummy1_send <= no_dummy1_send;
	no_dummy1_ack <= dummy1_ack;
	no_dummy1_rdy <= dummy1_rdy;
	dummy1_count <= no_dummy1_count;
	dummy2_data <= no_dummy2_data;
	dummy2_send <= no_dummy2_send;
	no_dummy2_ack <= dummy2_ack;
	no_dummy2_rdy <= dummy2_rdy;
	dummy2_count <= no_dummy2_count;
	dummy3_data <= no_dummy3_data;
	dummy3_send <= no_dummy3_send;
	no_dummy3_ack <= dummy3_ack;
	no_dummy3_rdy <= dummy3_rdy;
	dummy3_count <= no_dummy3_count;
	dummy4_data <= no_dummy4_data;
	dummy4_send <= no_dummy4_send;
	no_dummy4_ack <= dummy4_ack;
	no_dummy4_rdy <= dummy4_rdy;
	dummy4_count <= no_dummy4_count;
	
	-- Input Port(s) Instantiation
	ni_In_data <= In_data;
	ni_In_send <= In_send;
	In_ack <= ni_In_ack;
	In_rdy <= ni_In_rdy;
	ni_In_count <= In_count;
end architecture rtl;
-- ----------------------------------------------------------------------------
-- ----------------------------------------------------------------------------
-- ----------------------------------------------------------------------------
