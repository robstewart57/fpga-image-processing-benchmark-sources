// __  ___ __ ___  _ __   ___  ___ 
// \ \/ / '__/ _ \| '_ \ / _ \/ __|
//  >  <| | | (_) | | | | (_) \__ \
// /_/\_\_|  \___/|_| |_|\___/|___/
// 
// Xronos synthesizer version
// Run date: Thu 2 Nov 2017 13:57:13 +0000
// 

module LL1_L_iunzipFilter2D(Out2_COUNT, Out2_ACK, Out1_SEND, Out1_ACK, Out1_RDY, Out1_DATA, Out1_COUNT, Out2_RDY, In1_DATA, In1_ACK, In1_COUNT, RESET, CLK, In1_SEND, Out2_SEND, Out2_DATA);
wire		topLeft_done;
output	[15:0]	Out2_COUNT;
wire		midLeftNoConsume2_go;
wire		bottomRightNoConsume1_go;
wire		bottomRowNoConsume1_go;
wire		bottomRowNoConsume2_done;
wire		bottomLeftNoConsume2_go;
wire		donePopulateBuffer_done;
wire		bottomLeftNoConsume1_go;
wire		bottomLeftNoConsume1_done;
wire		midLeft1_done;
wire		midLeftNoConsume2_done;
wire		midRightNoConsume1_go;
wire		midNoConsume1_done;
wire		topRight_go;
input		Out2_ACK;
wire		midRight2_go;
output		Out1_SEND;
input		Out1_ACK;
wire		bottomRightNoConsume2_done;
wire		midLeft2_go;
wire		midRight1_go;
wire		bottomRowNoConsume1_done;
input		Out1_RDY;
wire		midRightNoConsume2_done;
output	[15:0]	Out1_DATA;
wire		midLeft2_done;
output	[15:0]	Out1_COUNT;
wire		bottomRowNoConsume2_go;
wire		populateBuffer_go;
input		Out2_RDY;
wire		mid1_go;
wire		topLeft_go;
wire		bottomLeftNoConsume2_done;
wire		midRight2_done;
wire		mid1_done;
wire		midRight1_done;
wire		donePopulateBuffer_go;
input	[15:0]	In1_DATA;
output		In1_ACK;
input	[15:0]	In1_COUNT;
wire		topRow_go;
input		RESET;
wire		midRightNoConsume1_done;
wire		populateBuffer_done;
wire		topRight_done;
input		CLK;
wire		mid2_done;
wire		midNoConsume1_go;
wire		midRightNoConsume2_go;
input		In1_SEND;
wire		topRow_done;
output		Out2_SEND;
wire		midLeftNoConsume1_go;
wire		mid2_go;
wire		midNoConsume2_done;
wire		bottomRightNoConsume2_go;
wire		bottomRightNoConsume1_done;
wire		midLeft1_go;
wire		midNoConsume2_go;
output	[15:0]	Out2_DATA;
wire		midLeftNoConsume1_done;
wire		bus_01bbf334_;
wire		scheduler_u59;
wire		scheduler_u67;
wire		scheduler_u60;
wire		LL1_L_iunzipFilter2D_scheduler_instance_DONE;
wire		scheduler_u56;
wire		scheduler_u55;
wire		scheduler_u74;
wire	[2:0]	scheduler_u54;
wire		scheduler_u57;
wire		scheduler_u65;
wire		scheduler_u66;
wire		scheduler;
wire		scheduler_u61;
wire		scheduler_u64;
wire		scheduler_u76;
wire		scheduler_u73;
wire		scheduler_u70;
wire		scheduler_u63;
wire		scheduler_u62;
wire		scheduler_u69;
wire		scheduler_u75;
wire		scheduler_u72;
wire		scheduler_u68;
wire		scheduler_u71;
wire		scheduler_u58;
wire		scheduler_u77;
wire		LL1_L_iunzipFilter2D_bottomLeftNoConsume1_instance_DONE;
wire		bottomLeftNoConsume1_u17;
wire		bottomLeftNoConsume1_u12;
wire		bottomLeftNoConsume1;
wire	[31:0]	bottomLeftNoConsume1_u13;
wire	[15:0]	bottomLeftNoConsume1_u11;
wire		bottomLeftNoConsume1_u10;
wire	[2:0]	bottomLeftNoConsume1_u14;
wire	[15:0]	bottomLeftNoConsume1_u9;
wire	[15:0]	bottomLeftNoConsume1_u16;
wire	[15:0]	bottomLeftNoConsume1_u15;
wire	[15:0]	bus_20897fac_;
wire		bus_0ca0f630_;
wire	[15:0]	bus_0ed5862c_;
wire		bus_1faaec31_;
wire	[15:0]	bus_4a9b702b_;
wire	[15:0]	bus_0cb909ae_;
wire	[15:0]	bus_3381d539_;
wire		bus_1ea2aac1_;
wire		bus_54485535_;
wire		bus_5858632d_;
wire	[15:0]	bus_47d6ef03_;
wire	[15:0]	bus_5f8b3986_;
wire	[15:0]	bus_232e245b_;
wire		bus_1ee56c59_;
wire		bus_349b9fac_;
wire		bus_6fff4e52_;
wire	[15:0]	bus_7351412b_;
wire	[15:0]	bus_694f6a4e_;
wire	[15:0]	bus_4c69ce54_;
wire	[15:0]	bus_55e3cbdb_;
wire		bus_12ab3e35_;
wire	[15:0]	bus_2ae9753e_;
wire	[15:0]	bus_01a2865d_;
wire	[15:0]	bus_06fef45c_;
wire	[15:0]	bus_28bb0475_;
wire		bus_1cb6406c_;
wire	[15:0]	bus_516e2378_;
wire		bus_013fe4a5_;
wire		bus_62557f73_;
wire		bus_59c5b7d5_;
wire	[15:0]	bus_42f56b99_;
wire		bus_600325c7_;
wire		bus_170909c9_;
wire		bus_34a996e5_;
wire	[15:0]	bus_3435fed4_;
wire		bus_05cc4bc4_;
wire		bus_18c7f89c_;
wire		bus_2bae7787_;
wire	[15:0]	bus_317adece_;
wire		bus_45e58a9c_;
wire	[31:0]	bus_1e0f9134_;
wire		bus_7f773641_;
wire		bus_3cc9da1f_;
wire		bus_5a2ebcef_;
wire	[15:0]	bus_7e595a89_;
wire	[15:0]	bus_4cbd1f1c_;
wire	[2:0]	bus_3607d9ee_;
wire		bus_6e4bea7e_;
wire		LL1_L_iunzipFilter2D_topRight_instance_DONE;
wire	[15:0]	topRight_u34;
wire	[15:0]	topRight_u24;
wire		topRight_u29;
wire		topRight_u27;
wire	[31:0]	topRight_u30;
wire		topRight;
wire	[2:0]	topRight_u35;
wire	[15:0]	topRight_u22;
wire	[15:0]	topRight_u37;
wire	[15:0]	topRight_u26;
wire	[31:0]	topRight_u33;
wire		topRight_u38;
wire		topRight_u28;
wire		topRight_u32;
wire		topRight_u23;
wire	[15:0]	topRight_u36;
wire		topRight_u39;
wire	[2:0]	topRight_u31;
wire		topRight_u21;
wire		topRight_u25;
wire	[31:0]	topRight_u20;
wire		bus_7290ab84_;
wire		or_6aa5e0aa_u0;
wire	[2:0]	midLeft2_u24;
wire	[15:0]	midLeft2_u30;
wire	[15:0]	midLeft2_u16;
wire		LL1_L_iunzipFilter2D_midLeft2_instance_DONE;
wire		midLeft2_u31;
wire		midLeft2_u19;
wire	[31:0]	midLeft2_u22;
wire		midLeft2_u29;
wire		midLeft2_u21;
wire		midLeft2;
wire	[31:0]	midLeft2_u26;
wire	[31:0]	midLeft2_u18;
wire		midLeft2_u25;
wire		midLeft2_u17;
wire	[15:0]	midLeft2_u28;
wire	[15:0]	midLeft2_u20;
wire	[15:0]	midLeft2_u23;
wire	[2:0]	midLeft2_u27;
wire	[15:0]	midLeftNoConsume2_u11;
wire	[31:0]	midLeftNoConsume2_u13;
wire		midLeftNoConsume2;
wire	[15:0]	midLeftNoConsume2_u9;
wire		midLeftNoConsume2_u12;
wire		midLeftNoConsume2_u16;
wire	[2:0]	midLeftNoConsume2_u14;
wire		midLeftNoConsume2_u10;
wire	[15:0]	midLeftNoConsume2_u17;
wire	[15:0]	midLeftNoConsume2_u15;
wire		LL1_L_iunzipFilter2D_midLeftNoConsume2_instance_DONE;
wire		bus_05b7360b_;
wire		bus_7ceb345f_;
wire		bottomLeftNoConsume2_u10;
wire		LL1_L_iunzipFilter2D_bottomLeftNoConsume2_instance_DONE;
wire		bottomLeftNoConsume2;
wire		bottomLeftNoConsume2_u12;
wire	[2:0]	bottomLeftNoConsume2_u14;
wire	[15:0]	bottomLeftNoConsume2_u11;
wire		bottomLeftNoConsume2_u17;
wire	[15:0]	bottomLeftNoConsume2_u9;
wire	[15:0]	bottomLeftNoConsume2_u15;
wire	[31:0]	bottomLeftNoConsume2_u13;
wire	[15:0]	bottomLeftNoConsume2_u16;
wire	[31:0]	topRow_u18;
wire	[15:0]	topRow_u20;
wire	[31:0]	topRow_u29;
wire	[15:0]	topRow_u32;
wire		LL1_L_iunzipFilter2D_topRow_instance_DONE;
wire		topRow_u25;
wire		topRow;
wire	[31:0]	topRow_u26;
wire		topRow_u23;
wire	[15:0]	topRow_u30;
wire		topRow_u19;
wire	[2:0]	topRow_u31;
wire	[15:0]	topRow_u24;
wire	[2:0]	topRow_u27;
wire		topRow_u28;
wire	[15:0]	topRow_u22;
wire	[15:0]	topRow_u33;
wire		topRow_u34;
wire		topRow_u21;
wire		topRow_u35;
wire		or_5aa0ea88_u0;
wire		bus_44ddb537_;
wire	[15:0]	bus_3ae80db9_;
wire		midRight1_u25;
wire	[15:0]	midRight1_u24;
wire	[31:0]	midRight1_u34;
wire	[31:0]	midRight1_u22;
wire		midRight1_u39;
wire	[15:0]	midRight1_u31;
wire		midRight1_u23;
wire		midRight1_u38;
wire		midRight1_u27;
wire	[15:0]	midRight1_u20;
wire	[15:0]	midRight1_u36;
wire		midRight1_u33;
wire		midRight1_u21;
wire	[2:0]	midRight1_u35;
wire		midRight1;
wire	[15:0]	midRight1_u37;
wire	[31:0]	midRight1_u30;
wire		midRight1_u29;
wire	[15:0]	midRight1_u26;
wire		midRight1_u28;
wire		LL1_L_iunzipFilter2D_midRight1_instance_DONE;
wire	[2:0]	midRight1_u32;
wire		bus_055a8fca_;
wire		bus_6b52f69a_;
wire		bus_434fd1c3_;
wire		bus_7fd1dd56_;
wire	[15:0]	midRight2_u20;
wire	[31:0]	midRight2_u22;
wire	[2:0]	midRight2_u35;
wire		midRight2_u25;
wire		midRight2;
wire	[15:0]	midRight2_u24;
wire	[31:0]	midRight2_u30;
wire		midRight2_u27;
wire	[15:0]	midRight2_u36;
wire		midRight2_u37;
wire	[15:0]	midRight2_u31;
wire		LL1_L_iunzipFilter2D_midRight2_instance_DONE;
wire	[2:0]	midRight2_u32;
wire		midRight2_u33;
wire		midRight2_u38;
wire	[15:0]	midRight2_u26;
wire		midRight2_u28;
wire	[31:0]	midRight2_u34;
wire		midRight2_u29;
wire	[15:0]	midRight2_u39;
wire		midRight2_u23;
wire		midRight2_u21;
wire	[15:0]	midLeft1_u16;
wire		midLeft1_u24;
wire	[15:0]	midLeft1_u20;
wire		midLeft1_u30;
wire		midLeft1_u19;
wire	[31:0]	midLeft1_u25;
wire		midLeft1_u21;
wire		midLeft1_u17;
wire		LL1_L_iunzipFilter2D_midLeft1_instance_DONE;
wire		midLeft1_u31;
wire	[2:0]	midLeft1_u27;
wire		midLeft1;
wire	[2:0]	midLeft1_u23;
wire	[15:0]	midLeft1_u26;
wire	[15:0]	midLeft1_u29;
wire	[31:0]	midLeft1_u22;
wire	[15:0]	midLeft1_u28;
wire	[31:0]	midLeft1_u18;
wire	[15:0]	bus_79ca6720_;
wire		bus_1e719960_;
wire		populateBuffer_u15;
wire		LL1_L_iunzipFilter2D_populateBuffer_instance_DONE;
wire		populateBuffer_u11;
wire		populateBuffer_u9;
wire	[15:0]	populateBuffer_u13;
wire	[31:0]	populateBuffer_u12;
wire	[15:0]	populateBuffer_u8;
wire	[31:0]	populateBuffer_u10;
wire		populateBuffer;
wire	[2:0]	populateBuffer_u14;
wire		mid1_u19;
wire		LL1_L_iunzipFilter2D_mid1_instance_DONE;
wire	[15:0]	mid1_u29;
wire	[31:0]	mid1_u22;
wire		mid1;
wire	[15:0]	mid1_u28;
wire		mid1_u17;
wire	[2:0]	mid1_u27;
wire		mid1_u24;
wire	[15:0]	mid1_u20;
wire		mid1_u30;
wire	[2:0]	mid1_u23;
wire	[15:0]	mid1_u18;
wire	[15:0]	mid1_u26;
wire	[31:0]	mid1_u16;
wire		mid1_u31;
wire		mid1_u21;
wire	[31:0]	mid1_u25;
wire		bus_36b55e90_;
wire		bus_55eeea99_;
wire		midNoConsume1_u12;
wire	[2:0]	midNoConsume1_u14;
wire	[31:0]	midNoConsume1_u13;
wire	[15:0]	midNoConsume1_u16;
wire	[15:0]	midNoConsume1_u9;
wire		midNoConsume1_u17;
wire		midNoConsume1_u10;
wire	[15:0]	midNoConsume1_u15;
wire		midNoConsume1;
wire		LL1_L_iunzipFilter2D_midNoConsume1_instance_DONE;
wire	[15:0]	midNoConsume1_u11;
wire		topLeft_u21;
wire		topLeft;
wire	[31:0]	topLeft_u18;
wire	[2:0]	topLeft_u23;
wire		topLeft_u30;
wire		topLeft_u19;
wire	[2:0]	topLeft_u27;
wire	[15:0]	topLeft_u29;
wire		topLeft_u31;
wire		topLeft_u24;
wire		LL1_L_iunzipFilter2D_topLeft_instance_DONE;
wire	[31:0]	topLeft_u22;
wire	[31:0]	topLeft_u25;
wire	[15:0]	topLeft_u28;
wire	[15:0]	topLeft_u16;
wire		topLeft_u17;
wire	[15:0]	topLeft_u26;
wire	[15:0]	topLeft_u20;
wire		donePopulateBuffer;
wire	[15:0]	donePopulateBuffer_u1;
wire		LL1_L_iunzipFilter2D_donePopulateBuffer_instance_DONE;
wire		bus_5a63b98e_;
wire		LL1_L_iunzipFilter2D_bottomRightNoConsume1_instance_DONE;
wire		bottomRightNoConsume1_u18;
wire	[15:0]	bottomRightNoConsume1_u17;
wire	[15:0]	bottomRightNoConsume1_u28;
wire		bottomRightNoConsume1_u20;
wire	[31:0]	bottomRightNoConsume1_u21;
wire	[15:0]	bottomRightNoConsume1_u27;
wire		bottomRightNoConsume1_u16;
wire		bottomRightNoConsume1;
wire		bottomRightNoConsume1_u23;
wire	[15:0]	bottomRightNoConsume1_u19;
wire		bottomRightNoConsume1_u24;
wire	[31:0]	bottomRightNoConsume1_u25;
wire	[2:0]	bottomRightNoConsume1_u26;
wire	[15:0]	bottomRightNoConsume1_u15;
wire		bottomRightNoConsume1_u29;
wire		bottomRightNoConsume1_u22;
wire		mid2_u31;
wire	[15:0]	mid2_u18;
wire	[31:0]	mid2_u25;
wire	[31:0]	mid2_u22;
wire		mid2_u29;
wire		mid2;
wire	[2:0]	mid2_u23;
wire		mid2_u17;
wire	[15:0]	mid2_u20;
wire		mid2_u24;
wire		mid2_u21;
wire	[15:0]	mid2_u26;
wire	[15:0]	mid2_u28;
wire		LL1_L_iunzipFilter2D_mid2_instance_DONE;
wire	[2:0]	mid2_u27;
wire	[15:0]	mid2_u30;
wire	[31:0]	mid2_u16;
wire		mid2_u19;
wire		midRightNoConsume1_u16;
wire		midRightNoConsume1;
wire		midRightNoConsume1_u15;
wire		LL1_L_iunzipFilter2D_midRightNoConsume1_instance_DONE;
wire	[15:0]	midRightNoConsume1_u13;
wire	[15:0]	midRightNoConsume1_u20;
wire		midRightNoConsume1_u21;
wire	[2:0]	midRightNoConsume1_u18;
wire	[31:0]	midRightNoConsume1_u17;
wire		midRightNoConsume1_u12;
wire	[15:0]	midRightNoConsume1_u19;
wire	[15:0]	midRightNoConsume1_u11;
wire		midRightNoConsume1_u14;
wire	[15:0]	bottomRowNoConsume1_u15;
wire	[15:0]	bottomRowNoConsume1_u9;
wire	[31:0]	bottomRowNoConsume1_u13;
wire		bottomRowNoConsume1_u10;
wire	[15:0]	bottomRowNoConsume1_u11;
wire		bottomRowNoConsume1;
wire		LL1_L_iunzipFilter2D_bottomRowNoConsume1_instance_DONE;
wire	[15:0]	bottomRowNoConsume1_u16;
wire		bottomRowNoConsume1_u17;
wire		bottomRowNoConsume1_u12;
wire	[2:0]	bottomRowNoConsume1_u14;
wire		bus_1e59a7e8_;
wire	[15:0]	bus_123b1c5f_;
wire		bus_33af7415_;
wire		bus_58ff9411_;
wire		bus_62c5dd82_;
wire	[2:0]	bus_31fab083_;
wire	[31:0]	bus_4b4b39e6_;
wire	[15:0]	or_0ed22344_u0;
wire		bus_74cef7bd_;
wire		bus_6e55ab9d_;
wire	[2:0]	bottomRowNoConsume2_u14;
wire	[15:0]	bottomRowNoConsume2_u11;
wire	[31:0]	bottomRowNoConsume2_u13;
wire		LL1_L_iunzipFilter2D_bottomRowNoConsume2_instance_DONE;
wire		bottomRowNoConsume2_u12;
wire	[15:0]	bottomRowNoConsume2_u9;
wire		bottomRowNoConsume2_u10;
wire	[15:0]	bottomRowNoConsume2_u15;
wire		bottomRowNoConsume2_u16;
wire	[15:0]	bottomRowNoConsume2_u17;
wire		bottomRowNoConsume2;
wire		bus_57d538ab_;
wire		bus_0e6b179e_;
wire		bus_4638b125_;
wire	[15:0]	bus_75e069b0_;
wire		bus_3e990c66_;
wire	[15:0]	bus_0189de6b_;
wire		bus_44ef805d_;
wire		bus_197870e1_;
wire		bus_4dd9231f_;
wire		bottomRightNoConsume2_u22;
wire		bottomRightNoConsume2_u23;
wire		bottomRightNoConsume2_u28;
wire		LL1_L_iunzipFilter2D_bottomRightNoConsume2_instance_DONE;
wire	[15:0]	bottomRightNoConsume2_u15;
wire	[15:0]	bottomRightNoConsume2_u27;
wire	[31:0]	bottomRightNoConsume2_u25;
wire		bottomRightNoConsume2_u20;
wire		bottomRightNoConsume2_u18;
wire		bottomRightNoConsume2;
wire		bottomRightNoConsume2_u16;
wire	[15:0]	bottomRightNoConsume2_u19;
wire	[15:0]	bottomRightNoConsume2_u29;
wire		bottomRightNoConsume2_u24;
wire	[15:0]	bottomRightNoConsume2_u17;
wire	[2:0]	bottomRightNoConsume2_u26;
wire	[31:0]	bottomRightNoConsume2_u21;
wire	[15:0]	bus_7da5ce18_;
wire		bus_6c6f8035_;
wire	[15:0]	bus_7a4ea340_;
wire	[15:0]	or_3f6158b1_u0;
wire	[15:0]	midRightNoConsume2_u20;
wire	[15:0]	midRightNoConsume2_u19;
wire		midRightNoConsume2_u12;
wire		midRightNoConsume2_u14;
wire	[2:0]	midRightNoConsume2_u18;
wire		midRightNoConsume2_u21;
wire	[15:0]	midRightNoConsume2_u11;
wire		midRightNoConsume2;
wire		midRightNoConsume2_u16;
wire	[31:0]	midRightNoConsume2_u17;
wire		LL1_L_iunzipFilter2D_midRightNoConsume2_instance_DONE;
wire	[15:0]	midRightNoConsume2_u13;
wire		midRightNoConsume2_u15;
wire		bus_15a8a0f9_;
wire		or_6e0c85d4_u0;
wire	[31:0]	bus_3d462f24_;
wire		bus_1e4fc043_;
wire	[2:0]	bus_5db5252c_;
wire	[15:0]	or_434270a3_u0;
wire		bus_595a4e1e_;
wire		midLeftNoConsume1_u12;
wire	[15:0]	midLeftNoConsume1_u11;
wire	[15:0]	midLeftNoConsume1_u9;
wire	[31:0]	midLeftNoConsume1_u13;
wire		midLeftNoConsume1_u17;
wire	[2:0]	midLeftNoConsume1_u14;
wire		LL1_L_iunzipFilter2D_midLeftNoConsume1_instance_DONE;
wire		midLeftNoConsume1_u10;
wire	[15:0]	midLeftNoConsume1_u16;
wire		midLeftNoConsume1;
wire	[15:0]	midLeftNoConsume1_u15;
wire	[15:0]	or_104a84be_u0;
wire	[31:0]	midNoConsume2_u13;
wire		midNoConsume2;
wire	[2:0]	midNoConsume2_u14;
wire		midNoConsume2_u17;
wire		midNoConsume2_u12;
wire		LL1_L_iunzipFilter2D_midNoConsume2_instance_DONE;
wire		midNoConsume2_u10;
wire	[15:0]	midNoConsume2_u11;
wire	[15:0]	midNoConsume2_u15;
wire	[15:0]	midNoConsume2_u16;
wire	[15:0]	midNoConsume2_u9;
assign topLeft_done=bus_36b55e90_;
assign Out2_COUNT=or_104a84be_u0;
assign midLeftNoConsume2_go=scheduler_u66;
assign bottomRightNoConsume1_go=scheduler_u68;
assign bottomRowNoConsume1_go=scheduler_u74;
assign bottomRowNoConsume2_done=bus_595a4e1e_;
assign bottomLeftNoConsume2_go=scheduler_u58;
assign donePopulateBuffer_done=bus_44ddb537_;
assign bottomLeftNoConsume1_go=scheduler_u61;
assign bottomLeftNoConsume1_done=bus_15a8a0f9_;
assign midLeft1_done=bus_7fd1dd56_;
assign midLeftNoConsume2_done=bus_6c6f8035_;
assign midRightNoConsume1_go=scheduler_u64;
assign midNoConsume1_done=bus_1e4fc043_;
assign topRight_go=scheduler_u72;
assign midRight2_go=scheduler_u75;
assign Out1_SEND=or_6aa5e0aa_u0;
assign bottomRightNoConsume2_done=bus_7ceb345f_;
assign midLeft2_go=scheduler_u59;
assign midRight1_go=scheduler_u60;
assign bottomRowNoConsume1_done=bus_74cef7bd_;
assign midRightNoConsume2_done=bus_4638b125_;
assign Out1_DATA=or_434270a3_u0;
assign midLeft2_done=bus_05b7360b_;
assign Out1_COUNT=or_0ed22344_u0;
assign bottomRowNoConsume2_go=scheduler_u77;
assign populateBuffer_go=scheduler_u55;
assign mid1_go=scheduler_u67;
assign topLeft_go=scheduler_u73;
assign bottomLeftNoConsume2_done=bus_4dd9231f_;
assign midRight2_done=bus_01bbf334_;
assign mid1_done=bus_0e6b179e_;
assign midRight1_done=bus_55eeea99_;
assign donePopulateBuffer_go=scheduler_u63;
assign In1_ACK=or_5aa0ea88_u0;
assign topRow_go=scheduler_u65;
assign midRightNoConsume1_done=bus_197870e1_;
assign populateBuffer_done=bus_6e55ab9d_;
assign topRight_done=bus_6e4bea7e_;
assign mid2_done=bus_5a63b98e_;
assign midNoConsume1_go=scheduler_u56;
assign midRightNoConsume2_go=scheduler_u57;
assign topRow_done=bus_57d538ab_;
assign Out2_SEND=or_6e0c85d4_u0;
assign midLeftNoConsume1_go=scheduler_u70;
assign mid2_go=scheduler_u76;
assign midNoConsume2_done=bus_1e719960_;
assign bottomRightNoConsume2_go=scheduler_u62;
assign bottomRightNoConsume1_done=bus_055a8fca_;
assign midLeft1_go=scheduler_u69;
assign midNoConsume2_go=scheduler_u71;
assign Out2_DATA=or_3f6158b1_u0;
assign midLeftNoConsume1_done=bus_434fd1c3_;
assign bus_01bbf334_=LL1_L_iunzipFilter2D_midRight2_instance_DONE&{1{LL1_L_iunzipFilter2D_midRight2_instance_DONE}};
LL1_L_iunzipFilter2D_scheduler LL1_L_iunzipFilter2D_scheduler_instance(.CLK(CLK), 
  .RESET(bus_7290ab84_), .GO(bus_1e59a7e8_), .port_2fdf62fc_(bus_5db5252c_), .port_3194e347_(bus_3ae80db9_), 
  .port_77e210a8_(bus_7da5ce18_), .port_1a03f6bd_(bus_7a4ea340_), .port_1d57b49c_(bus_3d462f24_), 
  .port_493b3a04_(bus_6b52f69a_), .port_4363ce38_(bottomRightNoConsume2_done), 
  .port_361addca_(In1_SEND), .port_3adbd198_(topLeft_done), .port_15705178_(midRight2_done), 
  .port_301c30b7_(topRow_done), .port_73f4be73_(mid1_done), .port_0d59c4af_(midRight1_done), 
  .port_79f2393c_(bottomRowNoConsume1_done), .port_687ecc25_(Out1_RDY), .port_37551257_(midRightNoConsume2_done), 
  .port_0a7c9fc4_(midLeft2_done), .port_7d10c806_(bottomRowNoConsume2_done), 
  .port_6cca95b7_(midNoConsume2_done), .port_30c305a6_(donePopulateBuffer_done), 
  .port_3f4943a6_(bottomLeftNoConsume1_done), .port_19c85cd4_(midLeft1_done), 
  .port_5b864c4b_(bottomRightNoConsume1_done), .port_4533a20c_(Out2_RDY), .port_39fe3b8f_(midLeftNoConsume2_done), 
  .port_4cf11580_(midNoConsume1_done), .port_4aa821f5_(midRightNoConsume1_done), 
  .port_4dced3ce_(populateBuffer_done), .port_56b37681_(bottomLeftNoConsume2_done), 
  .port_58e985b9_(topRight_done), .port_32814e4f_(midLeftNoConsume1_done), .port_56f644d1_(mid2_done), 
  .DONE(LL1_L_iunzipFilter2D_scheduler_instance_DONE), .RESULT(scheduler), .RESULT_u405(scheduler_u54), 
  .RESULT_u406(scheduler_u55), .RESULT_u407(scheduler_u56), .RESULT_u408(scheduler_u57), 
  .RESULT_u409(scheduler_u58), .RESULT_u410(scheduler_u59), .RESULT_u411(scheduler_u60), 
  .RESULT_u412(scheduler_u61), .RESULT_u413(scheduler_u62), .RESULT_u414(scheduler_u63), 
  .RESULT_u415(scheduler_u64), .RESULT_u416(scheduler_u65), .RESULT_u417(scheduler_u66), 
  .RESULT_u418(scheduler_u67), .RESULT_u419(scheduler_u68), .RESULT_u420(scheduler_u69), 
  .RESULT_u421(scheduler_u70), .RESULT_u422(scheduler_u71), .RESULT_u423(scheduler_u72), 
  .RESULT_u424(scheduler_u73), .RESULT_u425(scheduler_u74), .RESULT_u426(scheduler_u75), 
  .RESULT_u427(scheduler_u76), .RESULT_u428(scheduler_u77));
LL1_L_iunzipFilter2D_bottomLeftNoConsume1 LL1_L_iunzipFilter2D_bottomLeftNoConsume1_instance(.CLK(CLK), 
  .RESET(bus_7290ab84_), .GO(bottomLeftNoConsume1_go), .port_61b6f9d5_(16'h0), 
  .port_45192321_(bus_7da5ce18_), .port_068d9e17_(bus_6fff4e52_), .port_286032ff_(bus_0ed5862c_), 
  .DONE(LL1_L_iunzipFilter2D_bottomLeftNoConsume1_instance_DONE), .RESULT(bottomLeftNoConsume1), 
  .RESULT_u429(bottomLeftNoConsume1_u9), .RESULT_u430(bottomLeftNoConsume1_u10), 
  .RESULT_u431(bottomLeftNoConsume1_u11), .RESULT_u432(bottomLeftNoConsume1_u12), 
  .RESULT_u433(bottomLeftNoConsume1_u13), .RESULT_u434(bottomLeftNoConsume1_u14), 
  .RESULT_u435(bottomLeftNoConsume1_u15), .RESULT_u436(bottomLeftNoConsume1_u16), 
  .RESULT_u437(bottomLeftNoConsume1_u17));
LL1_L_iunzipFilter2D_simplememoryreferee_30774571_ LL1_L_iunzipFilter2D_simplememoryreferee_30774571__1(.bus_0243864e_(CLK), 
  .bus_5d3ae11e_(bus_7290ab84_), .bus_19484e64_(bus_3e990c66_), .bus_54e8abfe_(bus_75e069b0_), 
  .bus_20fb712d_(topLeft_u21), .bus_4f73f169_(topLeft_u24), .bus_4279a696_(topLeft_u26), 
  .bus_722d6b97_(topLeft_u25), .bus_1c777956_(3'h1), .bus_13f1caa2_(topRow_u25), 
  .bus_3bbec1a4_(topRow_u28), .bus_778a83e5_(topRow_u30), .bus_21b0d60f_(32'h0), 
  .bus_063abbd4_(3'h1), .bus_2b762ca1_(topRight_u29), .bus_5dfd93fb_(topRight_u32), 
  .bus_00516411_(topRight_u34), .bus_5370ed53_(32'h0), .bus_79564239_(3'h1), .bus_0e3a8226_(midLeft1_u21), 
  .bus_04a67cd7_(midLeft1_u24), .bus_460823b9_(midLeft1_u26), .bus_10bdbe2d_(32'h0), 
  .bus_4a03791e_(3'h1), .bus_51c5155e_(midLeft2_u25), .bus_23637f81_(midLeft2_u21), 
  .bus_23e6302d_(midLeft2_u23), .bus_6eb29e4f_(32'h0), .bus_613d1e04_(3'h1), .bus_5dcadfde_(midLeftNoConsume1_u12), 
  .bus_5c51a8d6_(32'h0), .bus_6767df53_(3'h1), .bus_6fa6325e_(midLeftNoConsume2_u12), 
  .bus_7167efe2_(32'h0), .bus_5884faca_(3'h1), .bus_7b82651c_(mid1_u21), .bus_12700c62_(mid1_u24), 
  .bus_78f2c71d_(mid1_u26), .bus_01cfc67d_(32'h0), .bus_69d0e5eb_(3'h1), .bus_3ae0aed4_(mid2_u21), 
  .bus_3f2f9d38_(mid2_u24), .bus_65a9722f_(mid2_u26), .bus_16b5d3be_(32'h0), .bus_45dfafc9_(3'h1), 
  .bus_35488083_(midNoConsume1_u12), .bus_7f794c6e_(32'h0), .bus_32e4169c_(3'h1), 
  .bus_7247ce17_(midNoConsume2_u12), .bus_3998d8b1_(32'h0), .bus_3df97d91_(3'h1), 
  .bus_5c6c776e_(midRight1_u33), .bus_5ab9a6be_(midRight1_u29), .bus_2d128350_(midRight1_u31), 
  .bus_54e5d40a_(32'h0), .bus_3246468e_(3'h1), .bus_4a5121f7_(midRight2_u33), .bus_5c683fe8_(midRight2_u29), 
  .bus_3189a35f_(midRight2_u31), .bus_1c1d4898_(32'h0), .bus_224fa6f5_(3'h1), .bus_6a39073c_(midRightNoConsume1_u16), 
  .bus_06490750_(32'h0), .bus_22f52c59_(3'h1), .bus_5ee61a28_(midRightNoConsume2_u16), 
  .bus_17b97c76_(32'h0), .bus_2346e771_(3'h1), .bus_21b39f31_(bottomLeftNoConsume1_u12), 
  .bus_15a2faf2_(32'h0), .bus_6ab9c209_(3'h1), .bus_59a547a4_(bottomLeftNoConsume2_u12), 
  .bus_2eda6c29_(32'h0), .bus_3121b847_(3'h1), .bus_75ed37c9_(bottomRowNoConsume1_u12), 
  .bus_7bb56cf6_(32'h0), .bus_577fde87_(3'h1), .bus_0b12336f_(bottomRowNoConsume2_u12), 
  .bus_711297cf_(32'h0), .bus_4a8a2bdd_(3'h1), .bus_5968c0b8_(bottomRightNoConsume1_u24), 
  .bus_15eaab9b_(32'h0), .bus_14b7951c_(3'h1), .bus_4ab46008_(bottomRightNoConsume2_u24), 
  .bus_2f560388_(32'h0), .bus_2e43f4db_(3'h1), .bus_47d6ef03_(bus_47d6ef03_), .bus_1e0f9134_(bus_1e0f9134_), 
  .bus_7f773641_(bus_7f773641_), .bus_349b9fac_(bus_349b9fac_), .bus_3607d9ee_(bus_3607d9ee_), 
  .bus_28bb0475_(bus_28bb0475_), .bus_170909c9_(bus_170909c9_), .bus_4c69ce54_(bus_4c69ce54_), 
  .bus_1ea2aac1_(bus_1ea2aac1_), .bus_20897fac_(bus_20897fac_), .bus_05cc4bc4_(bus_05cc4bc4_), 
  .bus_694f6a4e_(bus_694f6a4e_), .bus_3cc9da1f_(bus_3cc9da1f_), .bus_232e245b_(bus_232e245b_), 
  .bus_1cb6406c_(bus_1cb6406c_), .bus_7351412b_(bus_7351412b_), .bus_45e58a9c_(bus_45e58a9c_), 
  .bus_06fef45c_(bus_06fef45c_), .bus_1faaec31_(bus_1faaec31_), .bus_3381d539_(bus_3381d539_), 
  .bus_0ca0f630_(bus_0ca0f630_), .bus_317adece_(bus_317adece_), .bus_12ab3e35_(bus_12ab3e35_), 
  .bus_7e595a89_(bus_7e595a89_), .bus_18c7f89c_(bus_18c7f89c_), .bus_55e3cbdb_(bus_55e3cbdb_), 
  .bus_54485535_(bus_54485535_), .bus_4a9b702b_(bus_4a9b702b_), .bus_013fe4a5_(bus_013fe4a5_), 
  .bus_3435fed4_(bus_3435fed4_), .bus_1ee56c59_(bus_1ee56c59_), .bus_5f8b3986_(bus_5f8b3986_), 
  .bus_59c5b7d5_(bus_59c5b7d5_), .bus_2ae9753e_(bus_2ae9753e_), .bus_5a2ebcef_(bus_5a2ebcef_), 
  .bus_0ed5862c_(bus_0ed5862c_), .bus_6fff4e52_(bus_6fff4e52_), .bus_4cbd1f1c_(bus_4cbd1f1c_), 
  .bus_600325c7_(bus_600325c7_), .bus_0cb909ae_(bus_0cb909ae_), .bus_62557f73_(bus_62557f73_), 
  .bus_42f56b99_(bus_42f56b99_), .bus_2bae7787_(bus_2bae7787_), .bus_01a2865d_(bus_01a2865d_), 
  .bus_5858632d_(bus_5858632d_), .bus_516e2378_(bus_516e2378_), .bus_34a996e5_(bus_34a996e5_));
assign bus_6e4bea7e_=LL1_L_iunzipFilter2D_topRight_instance_DONE&{1{LL1_L_iunzipFilter2D_topRight_instance_DONE}};
LL1_L_iunzipFilter2D_topRight LL1_L_iunzipFilter2D_topRight_instance(.CLK(CLK), 
  .RESET(bus_7290ab84_), .GO(topRight_go), .port_441cd972_(bus_3d462f24_), .port_7fcde167_(bus_6b52f69a_), 
  .port_05ea2457_(bus_05cc4bc4_), .port_6215fb35_(bus_20897fac_), .port_4a4dafea_(bus_05cc4bc4_), 
  .port_50ff8e8d_(In1_DATA), .DONE(LL1_L_iunzipFilter2D_topRight_instance_DONE), 
  .RESULT(topRight), .RESULT_u438(topRight_u20), .RESULT_u439(topRight_u21), .RESULT_u440(topRight_u22), 
  .RESULT_u441(topRight_u23), .RESULT_u442(topRight_u24), .RESULT_u443(topRight_u25), 
  .RESULT_u444(topRight_u26), .RESULT_u445(topRight_u27), .RESULT_u446(topRight_u28), 
  .RESULT_u447(topRight_u29), .RESULT_u448(topRight_u30), .RESULT_u449(topRight_u31), 
  .RESULT_u450(topRight_u32), .RESULT_u451(topRight_u33), .RESULT_u452(topRight_u34), 
  .RESULT_u453(topRight_u35), .RESULT_u454(topRight_u36), .RESULT_u455(topRight_u37), 
  .RESULT_u456(topRight_u38), .RESULT_u457(topRight_u39));
LL1_L_iunzipFilter2D_globalreset_physical_3810141d_ LL1_L_iunzipFilter2D_globalreset_physical_3810141d__1(.bus_3dc23f78_(CLK), 
  .bus_2f4fdc33_(RESET), .bus_7290ab84_(bus_7290ab84_));
assign or_6aa5e0aa_u0=topLeft_u31|topRow_u35|topRight_u39|midLeft1_u31|midLeftNoConsume1_u17|mid1_u31|midNoConsume1_u17|midRight1_u39|midRightNoConsume1_u21|bottomLeftNoConsume1_u17|bottomRowNoConsume1_u17|bottomRightNoConsume1_u29;
LL1_L_iunzipFilter2D_midLeft2 LL1_L_iunzipFilter2D_midLeft2_instance(.CLK(CLK), 
  .RESET(bus_7290ab84_), .GO(midLeft2_go), .port_38ad9985_(16'h0), .port_56487516_(bus_3d462f24_), 
  .port_17d61741_(bus_7da5ce18_), .port_58424af2_(bus_1cb6406c_), .port_0d7c2f45_(bus_1cb6406c_), 
  .port_43399a57_(bus_232e245b_), .port_541437a9_(In1_DATA), .DONE(LL1_L_iunzipFilter2D_midLeft2_instance_DONE), 
  .RESULT(midLeft2), .RESULT_u458(midLeft2_u16), .RESULT_u459(midLeft2_u17), .RESULT_u460(midLeft2_u18), 
  .RESULT_u461(midLeft2_u19), .RESULT_u462(midLeft2_u20), .RESULT_u466(midLeft2_u21), 
  .RESULT_u467(midLeft2_u22), .RESULT_u468(midLeft2_u23), .RESULT_u469(midLeft2_u24), 
  .RESULT_u463(midLeft2_u25), .RESULT_u464(midLeft2_u26), .RESULT_u465(midLeft2_u27), 
  .RESULT_u470(midLeft2_u28), .RESULT_u471(midLeft2_u29), .RESULT_u472(midLeft2_u30), 
  .RESULT_u473(midLeft2_u31));
LL1_L_iunzipFilter2D_midLeftNoConsume2 LL1_L_iunzipFilter2D_midLeftNoConsume2_instance(.CLK(CLK), 
  .RESET(bus_7290ab84_), .GO(midLeftNoConsume2_go), .port_056011bc_(16'h0), .port_535b0b03_(bus_7da5ce18_), 
  .port_383828d2_(bus_1faaec31_), .port_1ffe318b_(bus_06fef45c_), .DONE(LL1_L_iunzipFilter2D_midLeftNoConsume2_instance_DONE), 
  .RESULT(midLeftNoConsume2), .RESULT_u474(midLeftNoConsume2_u9), .RESULT_u475(midLeftNoConsume2_u10), 
  .RESULT_u476(midLeftNoConsume2_u11), .RESULT_u477(midLeftNoConsume2_u12), .RESULT_u478(midLeftNoConsume2_u13), 
  .RESULT_u479(midLeftNoConsume2_u14), .RESULT_u480(midLeftNoConsume2_u15), .RESULT_u481(midLeftNoConsume2_u16), 
  .RESULT_u482(midLeftNoConsume2_u17));
assign bus_05b7360b_=LL1_L_iunzipFilter2D_midLeft2_instance_DONE&{1{LL1_L_iunzipFilter2D_midLeft2_instance_DONE}};
assign bus_7ceb345f_=LL1_L_iunzipFilter2D_bottomRightNoConsume2_instance_DONE&{1{LL1_L_iunzipFilter2D_bottomRightNoConsume2_instance_DONE}};
LL1_L_iunzipFilter2D_bottomLeftNoConsume2 LL1_L_iunzipFilter2D_bottomLeftNoConsume2_instance(.CLK(CLK), 
  .RESET(bus_7290ab84_), .GO(bottomLeftNoConsume2_go), .port_14deb7ac_(16'h0), 
  .port_68ceecfc_(bus_7da5ce18_), .port_3f625033_(bus_600325c7_), .port_1c9ca6f6_(bus_4cbd1f1c_), 
  .DONE(LL1_L_iunzipFilter2D_bottomLeftNoConsume2_instance_DONE), .RESULT(bottomLeftNoConsume2), 
  .RESULT_u483(bottomLeftNoConsume2_u9), .RESULT_u484(bottomLeftNoConsume2_u10), 
  .RESULT_u485(bottomLeftNoConsume2_u11), .RESULT_u486(bottomLeftNoConsume2_u12), 
  .RESULT_u487(bottomLeftNoConsume2_u13), .RESULT_u488(bottomLeftNoConsume2_u14), 
  .RESULT_u489(bottomLeftNoConsume2_u15), .RESULT_u490(bottomLeftNoConsume2_u16), 
  .RESULT_u491(bottomLeftNoConsume2_u17));
LL1_L_iunzipFilter2D_topRow LL1_L_iunzipFilter2D_topRow_instance(.CLK(CLK), .RESET(bus_7290ab84_), 
  .GO(topRow_go), .port_47a9ee1b_(bus_3d462f24_), .port_6d5aabbe_(bus_7da5ce18_), 
  .port_1f199a95_(bus_7a4ea340_), .port_2297a1f9_(bus_1ea2aac1_), .port_7ad5e7a2_(bus_4c69ce54_), 
  .port_7f824f8f_(bus_1ea2aac1_), .port_63075f82_(In1_DATA), .DONE(LL1_L_iunzipFilter2D_topRow_instance_DONE), 
  .RESULT(topRow), .RESULT_u492(topRow_u18), .RESULT_u493(topRow_u19), .RESULT_u494(topRow_u20), 
  .RESULT_u495(topRow_u21), .RESULT_u496(topRow_u22), .RESULT_u497(topRow_u23), 
  .RESULT_u498(topRow_u24), .RESULT_u499(topRow_u25), .RESULT_u500(topRow_u26), 
  .RESULT_u501(topRow_u27), .RESULT_u502(topRow_u28), .RESULT_u503(topRow_u29), 
  .RESULT_u504(topRow_u30), .RESULT_u505(topRow_u31), .RESULT_u506(topRow_u32), 
  .RESULT_u507(topRow_u33), .RESULT_u508(topRow_u34), .RESULT_u509(topRow_u35));
assign or_5aa0ea88_u0=populateBuffer_u15|topLeft_u30|topRow_u34|topRight_u38|midLeft1_u30|midLeft2_u29|mid1_u30|mid2_u29|midRight1_u38|midRight2_u37;
assign bus_44ddb537_=LL1_L_iunzipFilter2D_donePopulateBuffer_instance_DONE&{1{LL1_L_iunzipFilter2D_donePopulateBuffer_instance_DONE}};
LL1_L_iunzipFilter2D_stateVar_populatePtr LL1_L_iunzipFilter2D_stateVar_populatePtr_1(.bus_4bd01fea_(CLK), 
  .bus_5e5c669f_(bus_7290ab84_), .bus_5000423d_(populateBuffer), .bus_2631ddf5_(populateBuffer_u8), 
  .bus_2160680b_(donePopulateBuffer), .bus_338c8ca8_(16'h0), .bus_3ae80db9_(bus_3ae80db9_));
LL1_L_iunzipFilter2D_midRight1 LL1_L_iunzipFilter2D_midRight1_instance(.CLK(CLK), 
  .RESET(bus_7290ab84_), .GO(midRight1_go), .port_5255d759_(bus_3d462f24_), .port_14c39ecd_(bus_7a4ea340_), 
  .port_282e491b_(bus_6b52f69a_), .port_2c10671c_(bus_013fe4a5_), .port_4c76bba0_(bus_013fe4a5_), 
  .port_631edf34_(bus_4a9b702b_), .port_07cc4909_(In1_DATA), .DONE(LL1_L_iunzipFilter2D_midRight1_instance_DONE), 
  .RESULT(midRight1), .RESULT_u510(midRight1_u20), .RESULT_u511(midRight1_u21), 
  .RESULT_u512(midRight1_u22), .RESULT_u513(midRight1_u23), .RESULT_u514(midRight1_u24), 
  .RESULT_u515(midRight1_u25), .RESULT_u516(midRight1_u26), .RESULT_u517(midRight1_u27), 
  .RESULT_u518(midRight1_u28), .RESULT_u522(midRight1_u29), .RESULT_u523(midRight1_u30), 
  .RESULT_u524(midRight1_u31), .RESULT_u525(midRight1_u32), .RESULT_u519(midRight1_u33), 
  .RESULT_u520(midRight1_u34), .RESULT_u521(midRight1_u35), .RESULT_u526(midRight1_u36), 
  .RESULT_u527(midRight1_u37), .RESULT_u528(midRight1_u38), .RESULT_u529(midRight1_u39));
assign bus_055a8fca_=LL1_L_iunzipFilter2D_bottomRightNoConsume1_instance_DONE&{1{LL1_L_iunzipFilter2D_bottomRightNoConsume1_instance_DONE}};
LL1_L_iunzipFilter2D_stateVar_isEven LL1_L_iunzipFilter2D_stateVar_isEven_1(.bus_1f3489ff_(CLK), 
  .bus_4d0fbe00_(bus_7290ab84_), .bus_7316061a_(topRight_u27), .bus_78994a42_(topRight_u28), 
  .bus_52631b34_(midRight1_u27), .bus_1823e66f_(midRight1_u28), .bus_743d02cc_(midRight2_u27), 
  .bus_0a184a25_(midRight2_u28), .bus_40103492_(midRightNoConsume1_u14), .bus_7b46d837_(midRightNoConsume1_u15), 
  .bus_5dc6e0f1_(midRightNoConsume2_u14), .bus_1c6f5c87_(midRightNoConsume2_u15), 
  .bus_75eeb741_(bottomRightNoConsume1_u22), .bus_6f55ec5d_(bottomRightNoConsume1_u23), 
  .bus_581ab06d_(bottomRightNoConsume2_u22), .bus_51887cdb_(bottomRightNoConsume2_u23), 
  .bus_6b52f69a_(bus_6b52f69a_));
assign bus_434fd1c3_=LL1_L_iunzipFilter2D_midLeftNoConsume1_instance_DONE&{1{LL1_L_iunzipFilter2D_midLeftNoConsume1_instance_DONE}};
assign bus_7fd1dd56_=LL1_L_iunzipFilter2D_midLeft1_instance_DONE&{1{LL1_L_iunzipFilter2D_midLeft1_instance_DONE}};
LL1_L_iunzipFilter2D_midRight2 LL1_L_iunzipFilter2D_midRight2_instance(.CLK(CLK), 
  .RESET(bus_7290ab84_), .GO(midRight2_go), .port_7204953c_(bus_3d462f24_), .port_1cd54e3f_(bus_7a4ea340_), 
  .port_2166078e_(bus_6b52f69a_), .port_2a04576f_(bus_1ee56c59_), .port_38854079_(bus_1ee56c59_), 
  .port_1fe65f07_(bus_3435fed4_), .port_6e163b29_(In1_DATA), .DONE(LL1_L_iunzipFilter2D_midRight2_instance_DONE), 
  .RESULT(midRight2), .RESULT_u530(midRight2_u20), .RESULT_u531(midRight2_u21), 
  .RESULT_u532(midRight2_u22), .RESULT_u533(midRight2_u23), .RESULT_u534(midRight2_u24), 
  .RESULT_u535(midRight2_u25), .RESULT_u536(midRight2_u26), .RESULT_u537(midRight2_u27), 
  .RESULT_u538(midRight2_u28), .RESULT_u542(midRight2_u29), .RESULT_u543(midRight2_u30), 
  .RESULT_u544(midRight2_u31), .RESULT_u545(midRight2_u32), .RESULT_u539(midRight2_u33), 
  .RESULT_u540(midRight2_u34), .RESULT_u541(midRight2_u35), .RESULT_u546(midRight2_u36), 
  .RESULT_u547(midRight2_u37), .RESULT_u548(midRight2_u38), .RESULT_u549(midRight2_u39));
LL1_L_iunzipFilter2D_midLeft1 LL1_L_iunzipFilter2D_midLeft1_instance(.CLK(CLK), 
  .RESET(bus_7290ab84_), .GO(midLeft1_go), .port_250e58ba_(16'h0), .port_6197b3d4_(bus_3d462f24_), 
  .port_43ef7bd5_(bus_7da5ce18_), .port_36b60040_(bus_3cc9da1f_), .port_78b91e36_(bus_694f6a4e_), 
  .port_5a4c347c_(bus_3cc9da1f_), .port_616f0feb_(In1_DATA), .DONE(LL1_L_iunzipFilter2D_midLeft1_instance_DONE), 
  .RESULT(midLeft1), .RESULT_u550(midLeft1_u16), .RESULT_u551(midLeft1_u17), .RESULT_u552(midLeft1_u18), 
  .RESULT_u553(midLeft1_u19), .RESULT_u554(midLeft1_u20), .RESULT_u555(midLeft1_u21), 
  .RESULT_u556(midLeft1_u22), .RESULT_u557(midLeft1_u23), .RESULT_u558(midLeft1_u24), 
  .RESULT_u559(midLeft1_u25), .RESULT_u560(midLeft1_u26), .RESULT_u561(midLeft1_u27), 
  .RESULT_u562(midLeft1_u28), .RESULT_u563(midLeft1_u29), .RESULT_u564(midLeft1_u30), 
  .RESULT_u565(midLeft1_u31));
LL1_L_iunzipFilter2D_stateVar_idx LL1_L_iunzipFilter2D_stateVar_idx_1(.bus_62860c78_(CLK), 
  .bus_744fb394_(bus_7290ab84_), .bus_55af70f4_(topLeft), .bus_0ec28381_(16'h0), 
  .bus_7a64655b_(topRow_u19), .bus_25e2c4f7_(16'h0), .bus_3c68edfe_(topRight_u21), 
  .bus_04039d41_(16'h0), .bus_6208d411_(midLeft1), .bus_6483ddbc_(16'h0), .bus_7f2a89e4_(midLeft2), 
  .bus_6cd25c20_(16'h0), .bus_2fe413a1_(midLeftNoConsume1), .bus_77a210b0_(16'h0), 
  .bus_2ad73ea4_(midLeftNoConsume2), .bus_3f7de95e_(16'h0), .bus_0387bc2f_(mid1_u17), 
  .bus_61448fc8_(16'h0), .bus_7b1a01ba_(mid2_u17), .bus_12d790ff_(16'h0), .bus_69a6a217_(midNoConsume1), 
  .bus_539c4f12_(16'h0), .bus_1e9c9e19_(midNoConsume2), .bus_4104bb04_(16'h0), 
  .bus_48c5d111_(midRight1), .bus_50263840_(16'h0), .bus_1b1b4f63_(midRight2), 
  .bus_3d8d462c_(16'h0), .bus_03c74654_(bottomLeftNoConsume1), .bus_4c32e0b1_(16'h0), 
  .bus_0420cb9d_(bottomLeftNoConsume2), .bus_0f0be065_(16'h0), .bus_563eebef_(bottomRowNoConsume1), 
  .bus_6fc1dd73_(16'h0), .bus_1fe6e51c_(bottomRowNoConsume2), .bus_09922e92_(16'h0), 
  .bus_2fd9f75a_(bottomRightNoConsume1_u16), .bus_153933ae_(16'h0), .bus_0b1e2e3f_(bottomRightNoConsume2_u16), 
  .bus_61c6e306_(16'h0), .bus_79ca6720_(bus_79ca6720_));
assign bus_1e719960_=LL1_L_iunzipFilter2D_midNoConsume2_instance_DONE&{1{LL1_L_iunzipFilter2D_midNoConsume2_instance_DONE}};
LL1_L_iunzipFilter2D_populateBuffer LL1_L_iunzipFilter2D_populateBuffer_instance(.CLK(CLK), 
  .RESET(bus_7290ab84_), .GO(populateBuffer_go), .port_74e37b91_(bus_3ae80db9_), 
  .port_241c8e45_(bus_3d462f24_), .port_58f1a46c_(bus_33af7415_), .port_1a2c8dcf_(In1_DATA), 
  .DONE(LL1_L_iunzipFilter2D_populateBuffer_instance_DONE), .RESULT(populateBuffer), 
  .RESULT_u566(populateBuffer_u8), .RESULT_u567(populateBuffer_u9), .RESULT_u568(populateBuffer_u10), 
  .RESULT_u569(populateBuffer_u11), .RESULT_u570(populateBuffer_u12), .RESULT_u571(populateBuffer_u13), 
  .RESULT_u572(populateBuffer_u14), .RESULT_u573(populateBuffer_u15));
LL1_L_iunzipFilter2D_mid1 LL1_L_iunzipFilter2D_mid1_instance(.CLK(CLK), .RESET(bus_7290ab84_), 
  .GO(mid1_go), .port_60e25201_(bus_3d462f24_), .port_4fa18e7c_(bus_7da5ce18_), 
  .port_14295d04_(bus_0ca0f630_), .port_1a5e1c20_(bus_3381d539_), .port_10388e5c_(bus_0ca0f630_), 
  .port_5ccf9322_(In1_DATA), .DONE(LL1_L_iunzipFilter2D_mid1_instance_DONE), 
  .RESULT(mid1), .RESULT_u574(mid1_u16), .RESULT_u575(mid1_u17), .RESULT_u576(mid1_u18), 
  .RESULT_u577(mid1_u19), .RESULT_u578(mid1_u20), .RESULT_u579(mid1_u21), .RESULT_u580(mid1_u22), 
  .RESULT_u581(mid1_u23), .RESULT_u582(mid1_u24), .RESULT_u583(mid1_u25), .RESULT_u584(mid1_u26), 
  .RESULT_u585(mid1_u27), .RESULT_u586(mid1_u28), .RESULT_u587(mid1_u29), .RESULT_u588(mid1_u30), 
  .RESULT_u589(mid1_u31));
assign bus_36b55e90_=LL1_L_iunzipFilter2D_topLeft_instance_DONE&{1{LL1_L_iunzipFilter2D_topLeft_instance_DONE}};
assign bus_55eeea99_=LL1_L_iunzipFilter2D_midRight1_instance_DONE&{1{LL1_L_iunzipFilter2D_midRight1_instance_DONE}};
LL1_L_iunzipFilter2D_midNoConsume1 LL1_L_iunzipFilter2D_midNoConsume1_instance(.CLK(CLK), 
  .RESET(bus_7290ab84_), .GO(midNoConsume1_go), .port_60826727_(bus_7da5ce18_), 
  .port_2cb31f5d_(bus_18c7f89c_), .port_09dd1a6b_(bus_7e595a89_), .DONE(LL1_L_iunzipFilter2D_midNoConsume1_instance_DONE), 
  .RESULT(midNoConsume1), .RESULT_u590(midNoConsume1_u9), .RESULT_u591(midNoConsume1_u10), 
  .RESULT_u592(midNoConsume1_u11), .RESULT_u593(midNoConsume1_u12), .RESULT_u594(midNoConsume1_u13), 
  .RESULT_u595(midNoConsume1_u14), .RESULT_u596(midNoConsume1_u15), .RESULT_u597(midNoConsume1_u16), 
  .RESULT_u598(midNoConsume1_u17));
LL1_L_iunzipFilter2D_topLeft LL1_L_iunzipFilter2D_topLeft_instance(.CLK(CLK), 
  .RESET(bus_7290ab84_), .GO(topLeft_go), .port_37621793_(16'h0), .port_327d2b21_(bus_3d462f24_), 
  .port_25f1e81f_(bus_7da5ce18_), .port_2475269b_(bus_170909c9_), .port_0b3965ec_(bus_28bb0475_), 
  .port_4341b031_(bus_170909c9_), .port_65941495_(In1_DATA), .DONE(LL1_L_iunzipFilter2D_topLeft_instance_DONE), 
  .RESULT(topLeft), .RESULT_u599(topLeft_u16), .RESULT_u600(topLeft_u17), .RESULT_u601(topLeft_u18), 
  .RESULT_u602(topLeft_u19), .RESULT_u603(topLeft_u20), .RESULT_u604(topLeft_u21), 
  .RESULT_u605(topLeft_u22), .RESULT_u606(topLeft_u23), .RESULT_u607(topLeft_u24), 
  .RESULT_u608(topLeft_u25), .RESULT_u609(topLeft_u26), .RESULT_u610(topLeft_u27), 
  .RESULT_u611(topLeft_u28), .RESULT_u612(topLeft_u29), .RESULT_u613(topLeft_u30), 
  .RESULT_u614(topLeft_u31));
LL1_L_iunzipFilter2D_donePopulateBuffer LL1_L_iunzipFilter2D_donePopulateBuffer_instance(.CLK(CLK), 
  .RESET(bus_7290ab84_), .GO(donePopulateBuffer_go), .DONE(LL1_L_iunzipFilter2D_donePopulateBuffer_instance_DONE), 
  .RESULT(donePopulateBuffer), .RESULT_u615(donePopulateBuffer_u1));
assign bus_5a63b98e_=LL1_L_iunzipFilter2D_mid2_instance_DONE&{1{LL1_L_iunzipFilter2D_mid2_instance_DONE}};
LL1_L_iunzipFilter2D_bottomRightNoConsume1 LL1_L_iunzipFilter2D_bottomRightNoConsume1_instance(.CLK(CLK), 
  .RESET(bus_7290ab84_), .GO(bottomRightNoConsume1_go), .port_1bf2f003_(bus_6b52f69a_), 
  .port_727877ba_(bus_5858632d_), .port_16605d60_(bus_01a2865d_), .DONE(LL1_L_iunzipFilter2D_bottomRightNoConsume1_instance_DONE), 
  .RESULT(bottomRightNoConsume1), .RESULT_u616(bottomRightNoConsume1_u15), .RESULT_u617(bottomRightNoConsume1_u16), 
  .RESULT_u618(bottomRightNoConsume1_u17), .RESULT_u619(bottomRightNoConsume1_u18), 
  .RESULT_u620(bottomRightNoConsume1_u19), .RESULT_u621(bottomRightNoConsume1_u20), 
  .RESULT_u622(bottomRightNoConsume1_u21), .RESULT_u623(bottomRightNoConsume1_u22), 
  .RESULT_u624(bottomRightNoConsume1_u23), .RESULT_u625(bottomRightNoConsume1_u24), 
  .RESULT_u626(bottomRightNoConsume1_u25), .RESULT_u627(bottomRightNoConsume1_u26), 
  .RESULT_u628(bottomRightNoConsume1_u27), .RESULT_u629(bottomRightNoConsume1_u28), 
  .RESULT_u630(bottomRightNoConsume1_u29));
LL1_L_iunzipFilter2D_mid2 LL1_L_iunzipFilter2D_mid2_instance(.CLK(CLK), .RESET(bus_7290ab84_), 
  .GO(mid2_go), .port_02e503c9_(bus_3d462f24_), .port_2ff1ab3b_(bus_7da5ce18_), 
  .port_26472692_(bus_12ab3e35_), .port_160d8dbf_(bus_317adece_), .port_4827c421_(bus_12ab3e35_), 
  .port_564f706b_(In1_DATA), .DONE(LL1_L_iunzipFilter2D_mid2_instance_DONE), 
  .RESULT(mid2), .RESULT_u631(mid2_u16), .RESULT_u632(mid2_u17), .RESULT_u633(mid2_u18), 
  .RESULT_u634(mid2_u19), .RESULT_u635(mid2_u20), .RESULT_u636(mid2_u21), .RESULT_u637(mid2_u22), 
  .RESULT_u638(mid2_u23), .RESULT_u639(mid2_u24), .RESULT_u640(mid2_u25), .RESULT_u641(mid2_u26), 
  .RESULT_u642(mid2_u27), .RESULT_u643(mid2_u28), .RESULT_u644(mid2_u29), .RESULT_u645(mid2_u30), 
  .RESULT_u646(mid2_u31));
LL1_L_iunzipFilter2D_midRightNoConsume1 LL1_L_iunzipFilter2D_midRightNoConsume1_instance(.CLK(CLK), 
  .RESET(bus_7290ab84_), .GO(midRightNoConsume1_go), .port_78715e37_(bus_7a4ea340_), 
  .port_157318c1_(bus_6b52f69a_), .port_7b7c41d3_(bus_59c5b7d5_), .port_260281da_(bus_5f8b3986_), 
  .DONE(LL1_L_iunzipFilter2D_midRightNoConsume1_instance_DONE), .RESULT(midRightNoConsume1), 
  .RESULT_u647(midRightNoConsume1_u11), .RESULT_u648(midRightNoConsume1_u12), 
  .RESULT_u649(midRightNoConsume1_u13), .RESULT_u650(midRightNoConsume1_u14), 
  .RESULT_u651(midRightNoConsume1_u15), .RESULT_u652(midRightNoConsume1_u16), 
  .RESULT_u653(midRightNoConsume1_u17), .RESULT_u654(midRightNoConsume1_u18), 
  .RESULT_u655(midRightNoConsume1_u19), .RESULT_u656(midRightNoConsume1_u20), 
  .RESULT_u657(midRightNoConsume1_u21));
LL1_L_iunzipFilter2D_bottomRowNoConsume1 LL1_L_iunzipFilter2D_bottomRowNoConsume1_instance(.CLK(CLK), 
  .RESET(bus_7290ab84_), .GO(bottomRowNoConsume1_go), .port_090c0601_(bus_7da5ce18_), 
  .port_2afc9e1d_(bus_62557f73_), .port_0baaff02_(bus_0cb909ae_), .DONE(LL1_L_iunzipFilter2D_bottomRowNoConsume1_instance_DONE), 
  .RESULT(bottomRowNoConsume1), .RESULT_u658(bottomRowNoConsume1_u9), .RESULT_u659(bottomRowNoConsume1_u10), 
  .RESULT_u660(bottomRowNoConsume1_u11), .RESULT_u661(bottomRowNoConsume1_u12), 
  .RESULT_u662(bottomRowNoConsume1_u13), .RESULT_u663(bottomRowNoConsume1_u14), 
  .RESULT_u664(bottomRowNoConsume1_u15), .RESULT_u665(bottomRowNoConsume1_u16), 
  .RESULT_u666(bottomRowNoConsume1_u17));
LL1_L_iunzipFilter2D_Kicker_15 LL1_L_iunzipFilter2D_Kicker_15_1(.CLK(CLK), .RESET(bus_7290ab84_), 
  .bus_1e59a7e8_(bus_1e59a7e8_));
LL1_L_iunzipFilter2D_simplememoryreferee_570ba99f_ LL1_L_iunzipFilter2D_simplememoryreferee_570ba99f__1(.bus_24dbf5d8_(CLK), 
  .bus_1e68ee92_(bus_7290ab84_), .bus_42b63aee_(bus_44ef805d_), .bus_4d929d8d_(bus_0189de6b_), 
  .bus_0dc704d1_(populateBuffer_u11), .bus_35b4734c_(populateBuffer_u13), .bus_3ff68fd8_(populateBuffer_u12), 
  .bus_2e8e26fe_(3'h1), .bus_123b1c5f_(bus_123b1c5f_), .bus_4b4b39e6_(bus_4b4b39e6_), 
  .bus_58ff9411_(bus_58ff9411_), .bus_62c5dd82_(bus_62c5dd82_), .bus_31fab083_(bus_31fab083_), 
  .bus_33af7415_(bus_33af7415_));
assign or_0ed22344_u0=topLeft_u29|topRow_u33|topRight_u37|midLeft1_u29|midLeftNoConsume1_u16|mid1_u29|midNoConsume1_u16|midRight1_u37|midRightNoConsume1_u20|bottomLeftNoConsume1_u16|bottomRowNoConsume1_u16|bottomRightNoConsume1_u28;
assign bus_74cef7bd_=LL1_L_iunzipFilter2D_bottomRowNoConsume1_instance_DONE&{1{LL1_L_iunzipFilter2D_bottomRowNoConsume1_instance_DONE}};
assign bus_6e55ab9d_=LL1_L_iunzipFilter2D_populateBuffer_instance_DONE&{1{LL1_L_iunzipFilter2D_populateBuffer_instance_DONE}};
LL1_L_iunzipFilter2D_bottomRowNoConsume2 LL1_L_iunzipFilter2D_bottomRowNoConsume2_instance(.CLK(CLK), 
  .RESET(bus_7290ab84_), .GO(bottomRowNoConsume2_go), .port_72d40a34_(bus_7da5ce18_), 
  .port_2dfef218_(bus_2bae7787_), .port_1cd6730f_(bus_42f56b99_), .DONE(LL1_L_iunzipFilter2D_bottomRowNoConsume2_instance_DONE), 
  .RESULT(bottomRowNoConsume2), .RESULT_u667(bottomRowNoConsume2_u9), .RESULT_u668(bottomRowNoConsume2_u10), 
  .RESULT_u669(bottomRowNoConsume2_u11), .RESULT_u670(bottomRowNoConsume2_u12), 
  .RESULT_u671(bottomRowNoConsume2_u13), .RESULT_u672(bottomRowNoConsume2_u14), 
  .RESULT_u673(bottomRowNoConsume2_u15), .RESULT_u674(bottomRowNoConsume2_u16), 
  .RESULT_u675(bottomRowNoConsume2_u17));
assign bus_57d538ab_=LL1_L_iunzipFilter2D_topRow_instance_DONE&{1{LL1_L_iunzipFilter2D_topRow_instance_DONE}};
assign bus_0e6b179e_=LL1_L_iunzipFilter2D_mid1_instance_DONE&{1{LL1_L_iunzipFilter2D_mid1_instance_DONE}};
assign bus_4638b125_=LL1_L_iunzipFilter2D_midRightNoConsume2_instance_DONE&{1{LL1_L_iunzipFilter2D_midRightNoConsume2_instance_DONE}};
LL1_L_iunzipFilter2D_structuralmemory_01e37556_ LL1_L_iunzipFilter2D_structuralmemory_01e37556__1(.CLK_u1(CLK), 
  .bus_5916951f_(bus_7290ab84_), .bus_7f082c33_(bus_4b4b39e6_), .bus_2219040d_(3'h1), 
  .bus_4d72aca4_(bus_62c5dd82_), .bus_6b921393_(bus_58ff9411_), .bus_1b1b36f0_(bus_123b1c5f_), 
  .bus_75697e3b_(bus_1e0f9134_), .bus_369fe81a_(3'h1), .bus_0986c750_(bus_349b9fac_), 
  .bus_339c133a_(bus_7f773641_), .bus_4db85e66_(bus_47d6ef03_), .bus_0189de6b_(bus_0189de6b_), 
  .bus_44ef805d_(bus_44ef805d_), .bus_75e069b0_(bus_75e069b0_), .bus_3e990c66_(bus_3e990c66_));
assign bus_197870e1_=LL1_L_iunzipFilter2D_midRightNoConsume1_instance_DONE&{1{LL1_L_iunzipFilter2D_midRightNoConsume1_instance_DONE}};
assign bus_4dd9231f_=LL1_L_iunzipFilter2D_bottomLeftNoConsume2_instance_DONE&{1{LL1_L_iunzipFilter2D_bottomLeftNoConsume2_instance_DONE}};
LL1_L_iunzipFilter2D_bottomRightNoConsume2 LL1_L_iunzipFilter2D_bottomRightNoConsume2_instance(.CLK(CLK), 
  .RESET(bus_7290ab84_), .GO(bottomRightNoConsume2_go), .port_6ecd2cdc_(bus_6b52f69a_), 
  .port_0eaeaa28_(bus_34a996e5_), .port_3ee0a27c_(bus_516e2378_), .DONE(LL1_L_iunzipFilter2D_bottomRightNoConsume2_instance_DONE), 
  .RESULT(bottomRightNoConsume2), .RESULT_u676(bottomRightNoConsume2_u15), .RESULT_u677(bottomRightNoConsume2_u16), 
  .RESULT_u678(bottomRightNoConsume2_u17), .RESULT_u679(bottomRightNoConsume2_u18), 
  .RESULT_u680(bottomRightNoConsume2_u19), .RESULT_u681(bottomRightNoConsume2_u20), 
  .RESULT_u682(bottomRightNoConsume2_u21), .RESULT_u683(bottomRightNoConsume2_u22), 
  .RESULT_u684(bottomRightNoConsume2_u23), .RESULT_u685(bottomRightNoConsume2_u24), 
  .RESULT_u686(bottomRightNoConsume2_u25), .RESULT_u687(bottomRightNoConsume2_u26), 
  .RESULT_u688(bottomRightNoConsume2_u27), .RESULT_u689(bottomRightNoConsume2_u28), 
  .RESULT_u690(bottomRightNoConsume2_u29));
LL1_L_iunzipFilter2D_stateVar_midPtr LL1_L_iunzipFilter2D_stateVar_midPtr_1(.bus_38bd42c5_(CLK), 
  .bus_00f33b37_(bus_7290ab84_), .bus_53c01961_(topLeft_u19), .bus_188a6b35_(topLeft_u20), 
  .bus_16d1222c_(topRow_u21), .bus_122af5f2_(topRow_u22), .bus_01f7a039_(topRight_u23), 
  .bus_0aba6433_(16'h0), .bus_698b642e_(midLeft1_u19), .bus_2bc2559e_(midLeft1_u20), 
  .bus_43c76f68_(midLeft2_u19), .bus_0903fe04_(midLeft2_u20), .bus_7e6c4fd8_(midLeftNoConsume1_u10), 
  .bus_7955a617_(midLeftNoConsume1_u11), .bus_2551f507_(midLeftNoConsume2_u10), 
  .bus_1a0acc16_(midLeftNoConsume2_u11), .bus_723ff3dc_(mid1_u19), .bus_2d47447b_(mid1_u20), 
  .bus_1ed9e97d_(mid2_u19), .bus_62513a6e_(mid2_u20), .bus_0a10bc57_(midNoConsume1_u10), 
  .bus_02599f9e_(midNoConsume1_u11), .bus_4f97ace6_(midNoConsume2_u10), .bus_6a732550_(midNoConsume2_u11), 
  .bus_0a1ca6cd_(midRight1_u25), .bus_1a147c05_(16'h0), .bus_7becdf00_(midRight2_u25), 
  .bus_5fec891a_(16'h0), .bus_1fdda57d_(midRightNoConsume1_u12), .bus_4b200500_(16'h0), 
  .bus_1826a746_(midRightNoConsume2_u12), .bus_5ce7e0b1_(16'h0), .bus_0b07ce99_(bottomLeftNoConsume1_u10), 
  .bus_58e8f3e2_(bottomLeftNoConsume1_u11), .bus_79009f57_(bottomLeftNoConsume2_u10), 
  .bus_1603d043_(bottomLeftNoConsume2_u11), .bus_10233de4_(bottomRowNoConsume1_u10), 
  .bus_4bb9035f_(bottomRowNoConsume1_u11), .bus_087b7bab_(bottomRowNoConsume2_u10), 
  .bus_4abfcc53_(bottomRowNoConsume2_u11), .bus_6d53b8af_(bottomRightNoConsume1_u18), 
  .bus_6c7eeb69_(16'h0), .bus_13e6efa8_(bottomRightNoConsume2_u18), .bus_6b6720f0_(16'h0), 
  .bus_7da5ce18_(bus_7da5ce18_));
assign bus_6c6f8035_=LL1_L_iunzipFilter2D_midLeftNoConsume2_instance_DONE&{1{LL1_L_iunzipFilter2D_midLeftNoConsume2_instance_DONE}};
LL1_L_iunzipFilter2D_stateVar_processedRows LL1_L_iunzipFilter2D_stateVar_processedRows_1(.bus_50f9a42f_(CLK), 
  .bus_2540158d_(bus_7290ab84_), .bus_029cd39d_(topRow_u23), .bus_3a105536_(topRow_u24), 
  .bus_3b123367_(topRight_u25), .bus_52a23a90_(16'h1), .bus_178131c8_(midRight1_u23), 
  .bus_25bedb97_(midRight1_u24), .bus_1305960f_(midRight2_u23), .bus_7e5a3b31_(midRight2_u24), 
  .bus_6ba6e043_(midRightNoConsume1), .bus_30eeb15a_(midRightNoConsume1_u11), 
  .bus_5d02476d_(midRightNoConsume2), .bus_137b120f_(midRightNoConsume2_u11), 
  .bus_0d79e859_(bottomRightNoConsume1), .bus_406a29e0_(16'h0), .bus_3f13ae55_(bottomRightNoConsume2), 
  .bus_707ce562_(16'h0), .bus_7a4ea340_(bus_7a4ea340_));
assign or_3f6158b1_u0=midLeft2_u28|midLeftNoConsume2_u15|mid2_u28|midNoConsume2_u15|midRight2_u36|midRightNoConsume2_u19|bottomLeftNoConsume2_u15|bottomRowNoConsume2_u15|bottomRightNoConsume2_u27;
LL1_L_iunzipFilter2D_midRightNoConsume2 LL1_L_iunzipFilter2D_midRightNoConsume2_instance(.CLK(CLK), 
  .RESET(bus_7290ab84_), .GO(midRightNoConsume2_go), .port_79bca4ff_(bus_7a4ea340_), 
  .port_2d1fccd3_(bus_6b52f69a_), .port_79275d09_(bus_5a2ebcef_), .port_5fb2661f_(bus_2ae9753e_), 
  .DONE(LL1_L_iunzipFilter2D_midRightNoConsume2_instance_DONE), .RESULT(midRightNoConsume2), 
  .RESULT_u691(midRightNoConsume2_u11), .RESULT_u692(midRightNoConsume2_u12), 
  .RESULT_u693(midRightNoConsume2_u13), .RESULT_u694(midRightNoConsume2_u14), 
  .RESULT_u695(midRightNoConsume2_u15), .RESULT_u696(midRightNoConsume2_u16), 
  .RESULT_u697(midRightNoConsume2_u17), .RESULT_u698(midRightNoConsume2_u18), 
  .RESULT_u699(midRightNoConsume2_u19), .RESULT_u700(midRightNoConsume2_u20), 
  .RESULT_u701(midRightNoConsume2_u21));
assign bus_15a8a0f9_=LL1_L_iunzipFilter2D_bottomLeftNoConsume1_instance_DONE&{1{LL1_L_iunzipFilter2D_bottomLeftNoConsume1_instance_DONE}};
assign or_6e0c85d4_u0=midLeft2_u31|midLeftNoConsume2_u16|mid2_u31|midNoConsume2_u17|midRight2_u38|midRightNoConsume2_u21|bottomLeftNoConsume2_u17|bottomRowNoConsume2_u16|bottomRightNoConsume2_u28;
LL1_L_iunzipFilter2D_stateVar_consumed LL1_L_iunzipFilter2D_stateVar_consumed_1(.bus_7424c935_(CLK), 
  .bus_1123d441_(bus_7290ab84_), .bus_3f16ffcc_(populateBuffer_u9), .bus_6227a442_(populateBuffer_u10), 
  .bus_7b8e9386_(topLeft_u17), .bus_067c086b_(topLeft_u18), .bus_0dde284b_(topRow), 
  .bus_07d88328_(topRow_u18), .bus_652ccf5e_(topRight), .bus_48c0b833_(topRight_u20), 
  .bus_3323d058_(midLeft1_u17), .bus_606ed600_(midLeft1_u18), .bus_48687f49_(midLeft2_u17), 
  .bus_64ad0da3_(midLeft2_u18), .bus_2c867b3c_(mid1), .bus_7aacda2c_(mid1_u16), 
  .bus_3c7f9dca_(mid2), .bus_56028ff8_(mid2_u16), .bus_4fdd9249_(midRight1_u21), 
  .bus_5dd8910a_(midRight1_u22), .bus_17ac4f32_(midRight2_u21), .bus_2ca297c8_(midRight2_u22), 
  .bus_6b11aeca_(bottomRightNoConsume1_u20), .bus_3e36f63b_(32'h0), .bus_4b2a5c22_(bottomRightNoConsume2_u20), 
  .bus_55ce97a1_(32'h0), .bus_3d462f24_(bus_3d462f24_));
assign bus_1e4fc043_=LL1_L_iunzipFilter2D_midNoConsume1_instance_DONE&{1{LL1_L_iunzipFilter2D_midNoConsume1_instance_DONE}};
LL1_L_iunzipFilter2D_stateVar_fsmState_LL1_L_iunzipFilter2D LL1_L_iunzipFilter2D_stateVar_fsmState_LL1_L_iunzipFilter2D_1(.bus_345dfb8f_(CLK), 
  .bus_61dd5bb3_(bus_7290ab84_), .bus_6854f934_(scheduler), .bus_38852323_(scheduler_u54), 
  .bus_5db5252c_(bus_5db5252c_));
assign or_434270a3_u0=topLeft_u28|topRow_u32|topRight_u36|midLeft1_u28|midLeftNoConsume1_u15|mid1_u28|midNoConsume1_u15|midRight1_u36|midRightNoConsume1_u19|bottomLeftNoConsume1_u15|bottomRowNoConsume1_u15|bottomRightNoConsume1_u27;
assign bus_595a4e1e_=LL1_L_iunzipFilter2D_bottomRowNoConsume2_instance_DONE&{1{LL1_L_iunzipFilter2D_bottomRowNoConsume2_instance_DONE}};
LL1_L_iunzipFilter2D_midLeftNoConsume1 LL1_L_iunzipFilter2D_midLeftNoConsume1_instance(.CLK(CLK), 
  .RESET(bus_7290ab84_), .GO(midLeftNoConsume1_go), .port_5a8739a4_(16'h0), .port_75d6138f_(bus_7da5ce18_), 
  .port_13e22dd9_(bus_45e58a9c_), .port_78b51d4c_(bus_7351412b_), .DONE(LL1_L_iunzipFilter2D_midLeftNoConsume1_instance_DONE), 
  .RESULT(midLeftNoConsume1), .RESULT_u702(midLeftNoConsume1_u9), .RESULT_u703(midLeftNoConsume1_u10), 
  .RESULT_u704(midLeftNoConsume1_u11), .RESULT_u705(midLeftNoConsume1_u12), .RESULT_u706(midLeftNoConsume1_u13), 
  .RESULT_u707(midLeftNoConsume1_u14), .RESULT_u708(midLeftNoConsume1_u15), .RESULT_u709(midLeftNoConsume1_u16), 
  .RESULT_u710(midLeftNoConsume1_u17));
assign or_104a84be_u0=midLeft2_u30|midLeftNoConsume2_u17|mid2_u30|midNoConsume2_u16|midRight2_u39|midRightNoConsume2_u20|bottomLeftNoConsume2_u16|bottomRowNoConsume2_u17|bottomRightNoConsume2_u29;
LL1_L_iunzipFilter2D_midNoConsume2 LL1_L_iunzipFilter2D_midNoConsume2_instance(.CLK(CLK), 
  .RESET(bus_7290ab84_), .GO(midNoConsume2_go), .port_0df859e8_(bus_7da5ce18_), 
  .port_3e58b459_(bus_54485535_), .port_14715090_(bus_55e3cbdb_), .DONE(LL1_L_iunzipFilter2D_midNoConsume2_instance_DONE), 
  .RESULT(midNoConsume2), .RESULT_u711(midNoConsume2_u9), .RESULT_u712(midNoConsume2_u10), 
  .RESULT_u713(midNoConsume2_u11), .RESULT_u714(midNoConsume2_u12), .RESULT_u715(midNoConsume2_u13), 
  .RESULT_u716(midNoConsume2_u14), .RESULT_u717(midNoConsume2_u15), .RESULT_u718(midNoConsume2_u16), 
  .RESULT_u719(midNoConsume2_u17));
endmodule



module LL1_L_iunzipFilter2D_scheduler(CLK, RESET, GO, port_2fdf62fc_, port_3194e347_, port_77e210a8_, port_1a03f6bd_, port_1d57b49c_, port_493b3a04_, port_4363ce38_, port_361addca_, port_3adbd198_, port_15705178_, port_301c30b7_, port_73f4be73_, port_0d59c4af_, port_79f2393c_, port_687ecc25_, port_37551257_, port_0a7c9fc4_, port_7d10c806_, port_6cca95b7_, port_30c305a6_, port_3f4943a6_, port_19c85cd4_, port_5b864c4b_, port_4533a20c_, port_39fe3b8f_, port_4cf11580_, port_4aa821f5_, port_4dced3ce_, port_56b37681_, port_58e985b9_, port_32814e4f_, port_56f644d1_, RESULT, RESULT_u405, RESULT_u406, RESULT_u407, RESULT_u408, RESULT_u409, RESULT_u410, RESULT_u411, RESULT_u412, RESULT_u413, RESULT_u414, RESULT_u415, RESULT_u416, RESULT_u417, RESULT_u418, RESULT_u419, RESULT_u420, RESULT_u421, RESULT_u422, RESULT_u423, RESULT_u424, RESULT_u425, RESULT_u426, RESULT_u427, RESULT_u428, DONE);
input		CLK;
input		RESET;
input		GO;
input	[2:0]	port_2fdf62fc_;
input	[15:0]	port_3194e347_;
input	[15:0]	port_77e210a8_;
input	[15:0]	port_1a03f6bd_;
input	[31:0]	port_1d57b49c_;
input		port_493b3a04_;
input		port_4363ce38_;
input		port_361addca_;
input		port_3adbd198_;
input		port_15705178_;
input		port_301c30b7_;
input		port_73f4be73_;
input		port_0d59c4af_;
input		port_79f2393c_;
input		port_687ecc25_;
input		port_37551257_;
input		port_0a7c9fc4_;
input		port_7d10c806_;
input		port_6cca95b7_;
input		port_30c305a6_;
input		port_3f4943a6_;
input		port_19c85cd4_;
input		port_5b864c4b_;
input		port_4533a20c_;
input		port_39fe3b8f_;
input		port_4cf11580_;
input		port_4aa821f5_;
input		port_4dced3ce_;
input		port_56b37681_;
input		port_58e985b9_;
input		port_32814e4f_;
input		port_56f644d1_;
output		RESULT;
output	[2:0]	RESULT_u405;
output		RESULT_u406;
output		RESULT_u407;
output		RESULT_u408;
output		RESULT_u409;
output		RESULT_u410;
output		RESULT_u411;
output		RESULT_u412;
output		RESULT_u413;
output		RESULT_u414;
output		RESULT_u415;
output		RESULT_u416;
output		RESULT_u417;
output		RESULT_u418;
output		RESULT_u419;
output		RESULT_u420;
output		RESULT_u421;
output		RESULT_u422;
output		RESULT_u423;
output		RESULT_u424;
output		RESULT_u425;
output		RESULT_u426;
output		RESULT_u427;
output		RESULT_u428;
output		DONE;
wire		and_u717_u0;
wire signed	[15:0]	lessThan_b_signed;
wire		lessThan;
wire signed	[15:0]	lessThan_a_signed;
wire signed	[15:0]	equals_b_signed;
wire		equals;
wire signed	[15:0]	equals_a_signed;
wire	[15:0]	lessThan_u19_a_unsigned;
wire	[15:0]	lessThan_u19_b_unsigned;
wire		lessThan_u19;
wire	[15:0]	equals_u40_a_unsigned;
wire		equals_u40;
wire	[15:0]	equals_u40_b_unsigned;
wire	[15:0]	equals_u41_b_unsigned;
wire	[15:0]	equals_u41_a_unsigned;
wire		equals_u41;
wire signed	[15:0]	lessThan_u20_b_signed;
wire signed	[15:0]	lessThan_u20_a_signed;
wire		lessThan_u20;
wire		andOp;
wire	[31:0]	lessThan_u21_b_unsigned;
wire		lessThan_u21;
wire	[31:0]	lessThan_u21_a_unsigned;
wire		andOp_u54;
wire		andOp_u55;
wire	[15:0]	equals_u42_a_unsigned;
wire	[15:0]	equals_u42_b_unsigned;
wire		equals_u42;
wire		lessThan_u22;
wire signed	[15:0]	lessThan_u22_a_signed;
wire signed	[15:0]	lessThan_u22_b_signed;
wire		andOp_u56;
wire	[31:0]	lessThan_u23_a_unsigned;
wire	[31:0]	lessThan_u23_b_unsigned;
wire		lessThan_u23;
wire		andOp_u57;
wire		not_u144;
wire		andOp_u58;
wire	[15:0]	equals_u43_a_unsigned;
wire		equals_u43;
wire	[15:0]	equals_u43_b_unsigned;
wire signed	[15:0]	lessThan_u24_b_signed;
wire		lessThan_u24;
wire signed	[15:0]	lessThan_u24_a_signed;
wire		andOp_u59;
wire	[31:0]	equals_u44_b_unsigned;
wire		equals_u44;
wire	[31:0]	equals_u44_a_unsigned;
wire		andOp_u60;
wire		andOp_u61;
wire		equals_u45;
wire	[15:0]	equals_u45_a_unsigned;
wire	[15:0]	equals_u45_b_unsigned;
wire signed	[15:0]	lessThan_u25_a_signed;
wire		lessThan_u25;
wire signed	[15:0]	lessThan_u25_b_signed;
wire		andOp_u62;
wire		equals_u46;
wire	[31:0]	equals_u46_b_unsigned;
wire	[31:0]	equals_u46_a_unsigned;
wire		andOp_u63;
wire		not_u145;
wire		andOp_u64;
wire	[15:0]	lessThan_u26_b_unsigned;
wire		lessThan_u26;
wire	[15:0]	lessThan_u26_a_unsigned;
wire signed	[15:0]	lessThan_u27_b_signed;
wire		lessThan_u27;
wire signed	[15:0]	lessThan_u27_a_signed;
wire		andOp_u65;
wire	[31:0]	lessThan_u28_a_unsigned;
wire	[31:0]	lessThan_u28_b_unsigned;
wire		lessThan_u28;
wire		andOp_u66;
wire		andOp_u67;
wire		lessThan_u29;
wire	[15:0]	lessThan_u29_b_unsigned;
wire	[15:0]	lessThan_u29_a_unsigned;
wire		lessThan_u30;
wire signed	[15:0]	lessThan_u30_a_signed;
wire signed	[15:0]	lessThan_u30_b_signed;
wire		andOp_u68;
wire		lessThan_u31;
wire	[31:0]	lessThan_u31_b_unsigned;
wire	[31:0]	lessThan_u31_a_unsigned;
wire		andOp_u69;
wire		not_u146;
wire		andOp_u70;
wire	[15:0]	lessThan_u32_b_unsigned;
wire	[15:0]	lessThan_u32_a_unsigned;
wire		lessThan_u32;
wire		equals_u47;
wire	[31:0]	equals_u47_a_unsigned;
wire	[31:0]	equals_u47_b_unsigned;
wire		andOp_u71;
wire		andOp_u72;
wire	[15:0]	lessThan_u33_a_unsigned;
wire		lessThan_u33;
wire	[15:0]	lessThan_u33_b_unsigned;
wire	[31:0]	equals_u48_b_unsigned;
wire		equals_u48;
wire	[31:0]	equals_u48_a_unsigned;
wire		andOp_u73;
wire		not_u147;
wire		andOp_u74;
wire	[15:0]	equals_u49_b_unsigned;
wire	[15:0]	equals_u49_a_unsigned;
wire		equals_u49;
wire	[31:0]	lessThan_u34_a_unsigned;
wire		lessThan_u34;
wire	[31:0]	lessThan_u34_b_unsigned;
wire		andOp_u75;
wire		andOp_u76;
wire	[15:0]	equals_u50_b_unsigned;
wire		equals_u50;
wire	[15:0]	equals_u50_a_unsigned;
wire	[31:0]	lessThan_u35_a_unsigned;
wire	[31:0]	lessThan_u35_b_unsigned;
wire		lessThan_u35;
wire		andOp_u77;
wire		not_u148;
wire		andOp_u78;
wire	[15:0]	equals_u51_a_unsigned;
wire	[15:0]	equals_u51_b_unsigned;
wire		equals_u51;
wire	[31:0]	equals_u52_b_unsigned;
wire	[31:0]	equals_u52_a_unsigned;
wire		equals_u52;
wire		andOp_u79;
wire		andOp_u80;
wire	[15:0]	equals_u53_b_unsigned;
wire		equals_u53;
wire	[15:0]	equals_u53_a_unsigned;
wire	[31:0]	equals_u54_a_unsigned;
wire	[31:0]	equals_u54_b_unsigned;
wire		equals_u54;
wire		andOp_u81;
wire		not_u149;
wire		andOp_u82;
wire	[15:0]	equals_u55_a_unsigned;
wire	[15:0]	equals_u55_b_unsigned;
wire		equals_u55;
wire signed	[15:0]	equals_u56_a_signed;
wire		equals_u56;
wire signed	[15:0]	equals_u56_b_signed;
wire		andOp_u83;
wire	[31:0]	equals_u57_a_unsigned;
wire	[31:0]	equals_u57_b_unsigned;
wire		equals_u57;
wire		andOp_u84;
wire		andOp_u85;
wire		equals_u58;
wire	[15:0]	equals_u58_a_unsigned;
wire	[15:0]	equals_u58_b_unsigned;
wire		equals_u59;
wire signed	[15:0]	equals_u59_a_signed;
wire signed	[15:0]	equals_u59_b_signed;
wire		andOp_u86;
wire	[31:0]	equals_u60_a_unsigned;
wire		equals_u60;
wire	[31:0]	equals_u60_b_unsigned;
wire		andOp_u87;
wire		not_u150;
wire		andOp_u88;
wire	[15:0]	lessThan_u36_b_unsigned;
wire		lessThan_u36;
wire	[15:0]	lessThan_u36_a_unsigned;
wire	[31:0]	equals_u61_a_unsigned;
wire	[31:0]	equals_u61_b_unsigned;
wire		equals_u61;
wire		andOp_u89;
wire		andOp_u90;
wire	[15:0]	lessThan_u37_a_unsigned;
wire		lessThan_u37;
wire	[15:0]	lessThan_u37_b_unsigned;
wire	[31:0]	equals_u62_b_unsigned;
wire	[31:0]	equals_u62_a_unsigned;
wire		equals_u62;
wire		andOp_u91;
wire		not_u151;
wire		andOp_u92;
wire		equals_u63;
wire	[15:0]	equals_u63_b_unsigned;
wire	[15:0]	equals_u63_a_unsigned;
wire	[31:0]	equals_u64_a_unsigned;
wire	[31:0]	equals_u64_b_unsigned;
wire		equals_u64;
wire		andOp_u93;
wire		andOp_u94;
wire		equals_u65;
wire	[15:0]	equals_u65_a_unsigned;
wire	[15:0]	equals_u65_b_unsigned;
wire		equals_u66;
wire	[31:0]	equals_u66_b_unsigned;
wire	[31:0]	equals_u66_a_unsigned;
wire		andOp_u95;
wire		not_u152;
wire		andOp_u96;
wire signed	[31:0]	equals_u67_b_signed;
wire		equals_u67;
wire signed	[31:0]	equals_u67_a_signed;
wire		and_u718_u0;
wire		not_u153_u0;
wire		and_u719_u0;
wire		andOp_u97;
wire		and_u720_u0;
wire		and_u721_u0;
wire		not_u154_u0;
wire		simplePinWrite;
wire		not_u155_u0;
wire		and_u722_u0;
wire		and_u723_u0;
wire		simplePinWrite_u123;
wire		and_u724_u0;
wire		and_u725_u0;
wire		or_u184_u0;
wire	[2:0]	mux_u44;
wire		and_u726_u0;
wire		and_u727_u0;
wire signed	[31:0]	equals_u68_a_signed;
wire signed	[31:0]	equals_u68_b_signed;
wire		equals_u68;
wire		not_u156_u0;
wire		and_u728_u0;
wire		and_u729_u0;
wire		not_u157_u0;
wire		and_u730_u0;
wire		and_u731_u0;
wire		and_u732_u0;
wire		and_u733_u0;
wire		not_u158_u0;
wire		simplePinWrite_u124;
wire		and_u734_u0;
reg		reg_59eedaaa_u0=1'h0;
reg		reg_27b4c651_u0=1'h0;
reg		and_delayed_u35=1'h0;
reg		reg_4a42b705_u0=1'h0;
reg		and_delayed_result_delayed_u3=1'h0;
reg		reg_6cac83a7_u0=1'h0;
wire		or_u185_u0;
reg		reg_4a42b705_result_delayed_u0=1'h0;
wire		and_u735_u0;
reg		reg_094d88c9_u0=1'h0;
wire		and_u736_u0;
wire		or_u186_u0;
wire		and_u737_u0;
wire		or_u187_u0;
wire		and_u738_u0;
wire		and_u739_u0;
reg		and_delayed_u36_u0=1'h0;
wire signed	[31:0]	equals_u69_b_signed;
wire		equals_u69;
wire signed	[31:0]	equals_u69_a_signed;
wire		and_u740_u0;
wire		not_u159_u0;
wire		and_u741_u0;
wire		andOp_u98;
wire		and_u742_u0;
wire		and_u743_u0;
wire		not_u160_u0;
wire		and_u744_u0;
wire		and_u745_u0;
wire		not_u161_u0;
wire		simplePinWrite_u125;
reg		reg_0b7664d7_u0=1'h0;
wire		and_u746_u0;
reg		reg_3ad7a739_u0=1'h0;
reg		reg_1bc19411_u0=1'h0;
wire		and_u747_u0;
reg		reg_3ad7a739_result_delayed_u0=1'h0;
reg		reg_1b0e6c79_u0=1'h0;
reg		and_delayed_u37_u0=1'h0;
wire		or_u188_u0;
reg		reg_0b7664d7_result_delayed_u0=1'h0;
wire		andOp_u99;
wire		not_u162_u0;
wire		and_u748_u0;
wire		and_u749_u0;
wire		and_u750_u0;
wire		not_u163_u0;
wire		and_u751_u0;
wire		simplePinWrite_u126;
reg		reg_25e2a223_u0=1'h0;
reg		reg_25e2a223_result_delayed_u0=1'h0;
wire		or_u189_u0;
reg		reg_6cb55ed9_u0=1'h0;
reg		reg_7132143c_u0=1'h0;
reg		reg_6cb55ed9_result_delayed_u0=1'h0;
wire		and_u752_u0;
reg		and_delayed_u38_u0=1'h0;
wire		and_u753_u0;
reg		and_delayed_u39_u0=1'h0;
wire		and_u754_u0;
wire		or_u190_u0;
wire		and_u755_u0;
reg		and_delayed_u40_u0=1'h0;
wire		and_u756_u0;
wire	[2:0]	mux_u45_u0;
wire		or_u191_u0;
wire		or_u192_u0;
wire		and_u757_u0;
reg		reg_43562f66_u0=1'h0;
wire		or_u193_u0;
wire		and_u758_u0;
wire		and_u759_u0;
wire signed	[31:0]	equals_u70_b_signed;
wire		equals_u70;
wire signed	[31:0]	equals_u70_a_signed;
wire		not_u164_u0;
wire		and_u760_u0;
wire		and_u761_u0;
wire		andOp_u100;
wire		not_u165_u0;
wire		and_u762_u0;
wire		and_u763_u0;
wire		and_u764_u0;
wire		and_u765_u0;
wire		not_u166_u0;
wire		simplePinWrite_u127;
wire		and_u766_u0;
reg		reg_6f936df5_u0=1'h0;
wire		or_u194_u0;
reg		reg_5373c17a_u0=1'h0;
reg		reg_5373c17a_result_delayed_u0=1'h0;
reg		and_delayed_u41_u0=1'h0;
reg		reg_6f936df5_result_delayed_u0=1'h0;
reg		reg_6f936df5_result_delayed_result_delayed_u0=1'h0;
wire		and_u767_u0;
reg		reg_6f936df5_result_delayed_result_delayed_result_delayed_u0=1'h0;
wire		andOp_u101;
wire		and_u768_u0;
wire		not_u167_u0;
wire		and_u769_u0;
wire		and_u770_u0;
wire		not_u168_u0;
wire		and_u771_u0;
wire		simplePinWrite_u128;
reg		reg_74073fe4_u0=1'h0;
wire		and_u772_u0;
reg		reg_0eaacf63_u0=1'h0;
wire		or_u195_u0;
reg		and_delayed_u42_u0=1'h0;
reg		reg_3acc3e9c_u0=1'h0;
reg		reg_24425050_u0=1'h0;
wire		and_u773_u0;
reg		and_delayed_result_delayed_u4_u0=1'h0;
reg		reg_0eaacf63_result_delayed_u0=1'h0;
wire		and_u774_u0;
wire		and_u775_u0;
wire		not_u169_u0;
wire		and_u776_u0;
wire		and_u777_u0;
wire		not_u170_u0;
wire		simplePinWrite_u129;
reg		reg_774e2f4e_u0=1'h0;
reg		reg_1efbe559_u0=1'h0;
reg		reg_376a948f_u0=1'h0;
wire		and_u778_u0;
reg		reg_4094683f_u0=1'h0;
reg		reg_774e2f4e_result_delayed_u0=1'h0;
wire		or_u196_u0;
wire		and_u779_u0;
reg		and_delayed_u43_u0=1'h0;
wire		and_u780_u0;
wire		and_u781_u0;
wire		not_u171_u0;
wire		and_u782_u0;
wire		and_u783_u0;
wire		not_u172_u0;
wire		simplePinWrite_u130;
wire		and_u784_u0;
reg		reg_549c7b3d_u0=1'h0;
reg		reg_3da7ac05_u0=1'h0;
wire		or_u197_u0;
reg		and_delayed_u44_u0=1'h0;
reg		reg_549c7b3d_result_delayed_u0=1'h0;
wire		and_u785_u0;
reg		reg_3da7ac05_result_delayed_u0=1'h0;
reg		reg_3da7ac05_result_delayed_result_delayed_u0=1'h0;
wire		and_u786_u0;
wire		or_u198_u0;
wire		and_u787_u0;
reg		and_delayed_u45_u0=1'h0;
wire		or_u199_u0;
wire		or_u200_u0;
wire		and_u788_u0;
wire		and_u789_u0;
wire		or_u201_u0;
wire		and_u790_u0;
wire		or_u202_u0;
wire		and_u791_u0;
wire		or_u203_u0;
wire		or_u204_u0;
wire		and_u792_u0;
wire		and_u793_u0;
wire		or_u205_u0;
wire		and_u794_u0;
reg		reg_05c7e893_u0=1'h0;
wire		and_u795_u0;
wire signed	[31:0]	equals_u71_b_signed;
wire signed	[31:0]	equals_u71_a_signed;
wire		equals_u71;
wire		and_u796_u0;
wire		not_u173_u0;
wire		and_u797_u0;
wire		andOp_u102;
wire		and_u798_u0;
wire		and_u799_u0;
wire		not_u174_u0;
wire		and_u800_u0;
wire		and_u801_u0;
wire		not_u175_u0;
wire		simplePinWrite_u131;
wire		or_u206_u0;
reg		reg_3226eb2c_u0=1'h0;
reg		reg_23c4568f_u0=1'h0;
reg		reg_74ec09a7_u0=1'h0;
wire		and_u802_u0;
wire		and_u803_u0;
reg		reg_23c4568f_result_delayed_u0=1'h0;
reg		reg_648fa1fc_u0=1'h0;
reg		and_delayed_u46_u0=1'h0;
reg		reg_3226eb2c_result_delayed_u0=1'h0;
wire		andOp_u103;
wire		not_u176_u0;
wire		and_u804_u0;
wire		and_u805_u0;
wire		and_u806_u0;
wire		not_u177_u0;
wire		and_u807_u0;
wire		simplePinWrite_u132;
reg		reg_4fea946b_u0=1'h0;
wire		and_u808_u0;
reg		reg_6e00556b_u0=1'h0;
wire		or_u207_u0;
reg		reg_6e00556b_result_delayed_u0=1'h0;
reg		reg_309dfcec_u0=1'h0;
reg		and_delayed_u47_u0=1'h0;
reg		reg_7b04c971_u0=1'h0;
wire		and_u809_u0;
reg		reg_4fea946b_result_delayed_u0=1'h0;
wire		not_u178_u0;
wire		and_u810_u0;
wire		and_u811_u0;
wire		not_u179_u0;
wire		and_u812_u0;
wire		and_u813_u0;
wire		simplePinWrite_u133;
reg		reg_7cdd073f_u0=1'h0;
reg		reg_01b946ba_u0=1'h0;
reg		reg_01b946ba_result_delayed_u0=1'h0;
wire		and_u814_u0;
reg		reg_526cf179_u0=1'h0;
wire		or_u208_u0;
reg		and_delayed_u48_u0=1'h0;
wire		and_u815_u0;
reg		reg_7cdd073f_result_delayed_u0=1'h0;
wire		and_u816_u0;
wire		not_u180_u0;
wire		and_u817_u0;
wire		and_u818_u0;
wire		and_u819_u0;
wire		not_u181_u0;
wire		simplePinWrite_u134;
reg		reg_49ca584b_u0=1'h0;
reg		reg_033b743f_u0=1'h0;
wire		and_u820_u0;
wire		or_u209_u0;
reg		and_delayed_u49_u0=1'h0;
wire		and_u821_u0;
reg		reg_033b743f_result_delayed_u0=1'h0;
reg		and_delayed_u50_u0=1'h0;
reg		reg_49ca584b_result_delayed_u0=1'h0;
wire		andOp_u104;
wire		and_u822_u0;
wire		and_u823_u0;
wire		not_u182_u0;
wire		not_u183_u0;
wire		and_u824_u0;
wire		and_u825_u0;
wire		simplePinWrite_u135;
reg		reg_38c345e9_u0=1'h0;
wire		and_u826_u0;
reg		reg_0d74457a_u0=1'h0;
wire		and_u827_u0;
reg		reg_2f356d21_u0=1'h0;
reg		and_delayed_u51_u0=1'h0;
wire		or_u210_u0;
reg		reg_38c345e9_result_delayed_u0=1'h0;
reg		reg_0d74457a_result_delayed_u0=1'h0;
reg		reg_0d74457a_result_delayed_result_delayed_u0=1'h0;
wire		andOp_u105;
wire		not_u184_u0;
wire		and_u828_u0;
wire		and_u829_u0;
wire		not_u185_u0;
wire		and_u830_u0;
wire		and_u831_u0;
wire		simplePinWrite_u136;
reg		reg_317cd17d_u0=1'h0;
reg		reg_002dc3a9_u0=1'h0;
wire		or_u211_u0;
reg		reg_71ed30e6_u0=1'h0;
wire		and_u832_u0;
wire		and_u833_u0;
reg		reg_624de640_u0=1'h0;
reg		reg_317cd17d_result_delayed_u0=1'h0;
reg		and_delayed_u52_u0=1'h0;
reg		reg_71ed30e6_result_delayed_u0=1'h0;
wire		and_u834_u0;
wire		not_u186_u0;
wire		and_u835_u0;
wire		and_u836_u0;
wire		not_u187_u0;
wire		and_u837_u0;
wire		simplePinWrite_u137;
reg		reg_63fb95d2_u0=1'h0;
wire		or_u212_u0;
reg		reg_398c8621_u0=1'h0;
reg		reg_63fb95d2_result_delayed_u0=1'h0;
reg		reg_63fb95d2_result_delayed_result_delayed_u0=1'h0;
reg		reg_4529a71b_u0=1'h0;
wire		and_u838_u0;
wire		and_u839_u0;
reg		and_delayed_u53_u0=1'h0;
wire		and_u840_u0;
wire		and_u841_u0;
wire		not_u188_u0;
wire		and_u842_u0;
wire		and_u843_u0;
wire		not_u189_u0;
wire		simplePinWrite_u138;
reg		reg_420f216e_u0=1'h0;
reg		reg_6e40f982_u0=1'h0;
reg		reg_2d931bb0_u0=1'h0;
reg		reg_15a02ae4_u0=1'h0;
reg		reg_3b71b3f6_u0=1'h0;
reg		reg_2d931bb0_result_delayed_u0=1'h0;
wire		or_u213_u0;
wire		and_u844_u0;
wire		and_u845_u0;
wire		and_u846_u0;
reg		and_delayed_u54_u0=1'h0;
wire		and_u847_u0;
wire		or_u214_u0;
wire		or_u215_u0;
wire		or_u216_u0;
wire		and_u848_u0;
wire		and_u849_u0;
wire		or_u217_u0;
wire		or_u218_u0;
wire		and_u850_u0;
wire		and_u851_u0;
wire		and_u852_u0;
wire		or_u219_u0;
wire		or_u220_u0;
wire		and_u853_u0;
wire		and_u854_u0;
wire		or_u221_u0;
wire	[2:0]	mux_u46_u0;
wire		or_u222_u0;
wire		and_u855_u0;
wire		or_u223_u0;
wire		and_u856_u0;
wire		and_u857_u0;
wire	[2:0]	mux_u47_u0;
wire		or_u224_u0;
wire		and_u858_u0;
wire		or_u225_u0;
wire		or_u226_u0;
wire	[2:0]	mux_u48_u0;
wire		and_u859_u0;
wire	[2:0]	mux_u49_u0;
wire		or_u227_u0;
wire		and_u860_u0;
wire		or_u228_u0;
wire		and_u861_u0;
wire		and_u862_u0;
reg		reg_17b91f93_u0=1'h0;
wire		or_u229_u0;
wire		and_u863_u0;
wire signed	[31:0]	equals_u72_b_signed;
wire		equals_u72;
wire signed	[31:0]	equals_u72_a_signed;
wire		and_u864_u0;
wire		not_u190_u0;
wire		and_u865_u0;
wire		andOp_u106;
wire		and_u866_u0;
wire		and_u867_u0;
wire		not_u191_u0;
wire		not_u192_u0;
wire		and_u868_u0;
wire		and_u869_u0;
wire		simplePinWrite_u139;
wire		and_u870_u0;
wire		and_u871_u0;
reg		reg_62867c89_u0=1'h0;
reg		and_delayed_u55_u0=1'h0;
reg		reg_342b0dff_u0=1'h0;
wire		or_u230_u0;
reg		reg_342b0dff_result_delayed_u0=1'h0;
reg		reg_62867c89_result_delayed_u0=1'h0;
reg		and_delayed_result_delayed_u5_u0=1'h0;
reg		and_delayed_u56_u0=1'h0;
wire		andOp_u107;
wire		not_u193_u0;
wire		and_u872_u0;
wire		and_u873_u0;
wire		and_u874_u0;
wire		and_u875_u0;
wire		not_u194_u0;
wire		simplePinWrite_u140;
reg		reg_5c254b63_u0=1'h0;
wire		and_u876_u0;
reg		reg_122ac30d_u0=1'h0;
reg		reg_4dcbcd47_u0=1'h0;
wire		and_u877_u0;
reg		reg_5c254b63_result_delayed_u0=1'h0;
reg		and_delayed_u57_u0=1'h0;
reg		reg_4dcbcd47_result_delayed_u0=1'h0;
wire		or_u231_u0;
reg		and_delayed_u58_u0=1'h0;
wire		not_u195_u0;
wire		and_u878_u0;
wire		and_u879_u0;
wire		and_u880_u0;
wire		and_u881_u0;
wire		not_u196_u0;
wire		simplePinWrite_u141;
reg		reg_4aef9f0e_u0=1'h0;
reg		reg_77e48187_u0=1'h0;
reg		reg_4aef9f0e_result_delayed_u0=1'h0;
wire		or_u232_u0;
reg		reg_307315fd_u0=1'h0;
reg		reg_307315fd_result_delayed_u0=1'h0;
reg		reg_4aef9f0e_result_delayed_result_delayed_u0=1'h0;
wire		and_u882_u0;
wire		and_u883_u0;
wire		and_u884_u0;
wire		not_u197_u0;
wire		and_u885_u0;
wire		and_u886_u0;
wire		and_u887_u0;
wire		not_u198_u0;
wire		simplePinWrite_u142;
reg		reg_7ee43ce2_u0=1'h0;
reg		reg_32619689_u0=1'h0;
reg		reg_5416fdbe_u0=1'h0;
wire		or_u233_u0;
reg		reg_32619689_result_delayed_u0=1'h0;
wire		and_u888_u0;
wire		and_u889_u0;
reg		reg_7ee43ce2_result_delayed_u0=1'h0;
reg		and_delayed_u59_u0=1'h0;
wire		not_u199_u0;
wire		and_u890_u0;
wire		and_u891_u0;
wire		and_u892_u0;
wire		and_u893_u0;
wire		not_u200_u0;
wire		simplePinWrite_u143;
reg		reg_7a4edfae_u0=1'h0;
reg		reg_25cc270d_u0=1'h0;
reg		reg_5b6f804b_u0=1'h0;
wire		and_u894_u0;
wire		and_u895_u0;
reg		and_delayed_u60_u0=1'h0;
wire		or_u234_u0;
reg		and_delayed_u61_u0=1'h0;
reg		and_delayed_result_delayed_u6_u0=1'h0;
wire		and_u896_u0;
wire		not_u201_u0;
wire		and_u897_u0;
wire		and_u898_u0;
wire		not_u202_u0;
wire		and_u899_u0;
wire		simplePinWrite_u144;
reg		reg_07a24aa2_u0=1'h0;
reg		reg_5887a60e_u0=1'h0;
reg		reg_0281fc6b_u0=1'h0;
reg		reg_0281fc6b_result_delayed_u0=1'h0;
reg		reg_07a24aa2_result_delayed_u0=1'h0;
reg		reg_09dc81cd_u0=1'h0;
wire		and_u900_u0;
wire		and_u901_u0;
wire		or_u235_u0;
wire		and_u902_u0;
wire		and_u903_u0;
wire		or_u236_u0;
reg		and_delayed_u62_u0=1'h0;
wire		and_u904_u0;
wire		or_u237_u0;
wire		and_u905_u0;
wire		or_u238_u0;
wire		and_u906_u0;
wire	[2:0]	mux_u50_u0;
wire		or_u239_u0;
wire		and_u907_u0;
wire		or_u240_u0;
wire		and_u908_u0;
wire		or_u241_u0;
wire		and_u909_u0;
wire	[2:0]	mux_u51_u0;
wire		or_u242_u0;
wire		and_u910_u0;
wire		and_u911_u0;
wire		or_u243_u0;
wire	[2:0]	mux_u52_u0;
wire		or_u244_u0;
wire		and_u912_u0;
wire		or_u245_u0;
wire	[2:0]	mux_u53_u0;
wire		or_u246_u0;
wire		and_u913_u0;
wire		or_u247_u0;
wire		and_u914_u0;
reg		and_delayed_u63_u0=1'h0;
wire		and_u915_u0;
wire signed	[31:0]	equals_u73_b_signed;
wire signed	[31:0]	equals_u73_a_signed;
wire		equals_u73;
wire		and_u916_u0;
wire		not_u203_u0;
wire		and_u917_u0;
wire		and_u918_u0;
wire		not_u204_u0;
wire		and_u919_u0;
wire		and_u920_u0;
wire		not_u205_u0;
wire		and_u921_u0;
wire		simplePinWrite_u145;
wire		and_u922_u0;
reg		reg_5938427c_u0=1'h0;
reg		reg_3a61ec86_u0=1'h0;
wire		and_u923_u0;
reg		and_delayed_u64_u0=1'h0;
reg		and_delayed_u65_u0=1'h0;
wire		or_u248_u0;
reg		reg_5938427c_result_delayed_u0=1'h0;
reg		reg_5938427c_result_delayed_result_delayed_u0=1'h0;
wire		and_u924_u0;
wire		and_u925_u0;
wire		not_u206_u0;
wire		not_u207_u0;
wire		and_u926_u0;
wire		and_u927_u0;
wire		simplePinWrite_u146;
wire		and_u928_u0;
wire		or_u249_u0;
reg		reg_0c3b0433_u0=1'h0;
reg		and_delayed_u66_u0=1'h0;
reg		reg_5a1c7caf_u0=1'h0;
reg		and_delayed_result_delayed_u7_u0=1'h0;
reg		reg_0c3b0433_result_delayed_u0=1'h0;
reg		reg_0c3b0433_result_delayed_result_delayed_u0=1'h0;
wire		and_u929_u0;
wire		not_u208_u0;
wire		and_u930_u0;
wire		and_u931_u0;
wire		and_u932_u0;
wire		and_u933_u0;
wire		not_u209_u0;
wire		simplePinWrite_u147;
wire		and_u934_u0;
reg		reg_3fb682df_u0=1'h0;
reg		reg_513f5af6_u0=1'h0;
wire		or_u250_u0;
reg		reg_0b0fac36_u0=1'h0;
wire		and_u935_u0;
reg		and_delayed_u67_u0=1'h0;
reg		reg_3fb682df_result_delayed_u0=1'h0;
reg		reg_513f5af6_result_delayed_u0=1'h0;
wire		and_u936_u0;
wire		not_u210_u0;
wire		and_u937_u0;
wire		and_u938_u0;
wire		and_u939_u0;
wire		not_u211_u0;
wire		simplePinWrite_u148;
reg		reg_4ecbafa0_u0=1'h0;
reg		reg_78c90025_u0=1'h0;
wire		and_u940_u0;
wire		and_u941_u0;
reg		and_delayed_u68_u0=1'h0;
reg		reg_46014afb_u0=1'h0;
reg		reg_4ecbafa0_result_delayed_u0=1'h0;
reg		and_delayed_u69_u0=1'h0;
wire		or_u251_u0;
wire		and_u942_u0;
reg		and_delayed_u70_u0=1'h0;
wire		or_u252_u0;
wire		and_u943_u0;
wire		and_u944_u0;
wire		or_u253_u0;
wire		or_u254_u0;
wire		and_u945_u0;
wire	[2:0]	mux_u54_u0;
wire		or_u255_u0;
wire		and_u946_u0;
wire		or_u256_u0;
wire		and_u947_u0;
wire		or_u257_u0;
wire		and_u948_u0;
wire	[2:0]	mux_u55_u0;
wire		or_u258_u0;
wire		and_u949_u0;
wire		and_u950_u0;
wire		or_u259_u0;
reg		reg_42f13385_u0=1'h0;
wire		and_u951_u0;
wire		midLeftNoConsume2_go_merge;
wire		midLeft2_go_merge;
wire		scoreboard_090d27ac_and;
reg		scoreboard_090d27ac_reg4=1'h0;
reg		scoreboard_090d27ac_reg0=1'h0;
reg		scoreboard_090d27ac_reg3=1'h0;
wire		scoreboard_090d27ac_resOr2;
wire		scoreboard_090d27ac_resOr0;
reg		scoreboard_090d27ac_reg5=1'h0;
wire		scoreboard_090d27ac_resOr3;
reg		scoreboard_090d27ac_reg2=1'h0;
wire		scoreboard_090d27ac_resOr4;
wire		scoreboard_090d27ac_resOr5;
reg		scoreboard_090d27ac_reg1=1'h0;
wire		scoreboard_090d27ac_resOr1;
wire		bus_07c053e2_;
wire		midLeft1_go_merge;
wire		midLeftNoConsume1_go_merge;
wire	[2:0]	mux_u56_u0;
wire		or_u260_u0;
wire		or_u261_u0;
reg		reg_12346cc9_u0=1'h0;
reg		reg_12346cc9_result_delayed_u0=1'h0;
wire	[2:0]	mux_u57_u0;
wire		or_u262_u0;
assign and_u717_u0=or_u261_u0&or_u261_u0;
assign lessThan_a_signed=port_3194e347_;
assign lessThan_b_signed=16'h103;
assign lessThan=lessThan_a_signed<lessThan_b_signed;
assign equals_a_signed=port_3194e347_;
assign equals_b_signed=16'h103;
assign equals=equals_a_signed==equals_b_signed;
assign lessThan_u19_a_unsigned=port_77e210a8_;
assign lessThan_u19_b_unsigned=16'hff;
assign lessThan_u19=lessThan_u19_a_unsigned<lessThan_u19_b_unsigned;
assign equals_u40_a_unsigned=port_77e210a8_;
assign equals_u40_b_unsigned=16'hff;
assign equals_u40=equals_u40_a_unsigned==equals_u40_b_unsigned;
assign equals_u41_a_unsigned=port_77e210a8_;
assign equals_u41_b_unsigned=16'h0;
assign equals_u41=equals_u41_a_unsigned==equals_u41_b_unsigned;
assign lessThan_u20_a_signed=port_1a03f6bd_;
assign lessThan_u20_b_signed=16'h1ff;
assign lessThan_u20=lessThan_u20_a_signed<lessThan_u20_b_signed;
assign andOp=equals_u41&lessThan_u20;
assign lessThan_u21_a_unsigned=port_1d57b49c_;
assign lessThan_u21_b_unsigned=32'h20000;
assign lessThan_u21=lessThan_u21_a_unsigned<lessThan_u21_b_unsigned;
assign andOp_u54=andOp&lessThan_u21;
assign andOp_u55=andOp_u54&port_493b3a04_;
assign equals_u42_a_unsigned=port_77e210a8_;
assign equals_u42_b_unsigned=16'h0;
assign equals_u42=equals_u42_a_unsigned==equals_u42_b_unsigned;
assign lessThan_u22_a_signed=port_1a03f6bd_;
assign lessThan_u22_b_signed=16'h1ff;
assign lessThan_u22=lessThan_u22_a_signed<lessThan_u22_b_signed;
assign andOp_u56=equals_u42&lessThan_u22;
assign lessThan_u23_a_unsigned=port_1d57b49c_;
assign lessThan_u23_b_unsigned=32'h20000;
assign lessThan_u23=lessThan_u23_a_unsigned<lessThan_u23_b_unsigned;
assign andOp_u57=andOp_u56&lessThan_u23;
assign not_u144=!port_493b3a04_;
assign andOp_u58=andOp_u57&not_u144;
assign equals_u43_a_unsigned=port_77e210a8_;
assign equals_u43_b_unsigned=16'h0;
assign equals_u43=equals_u43_a_unsigned==equals_u43_b_unsigned;
assign lessThan_u24_a_signed=port_1a03f6bd_;
assign lessThan_u24_b_signed=16'h1ff;
assign lessThan_u24=lessThan_u24_a_signed<lessThan_u24_b_signed;
assign andOp_u59=equals_u43&lessThan_u24;
assign equals_u44_a_unsigned=port_1d57b49c_;
assign equals_u44_b_unsigned=32'h20000;
assign equals_u44=equals_u44_a_unsigned==equals_u44_b_unsigned;
assign andOp_u60=andOp_u59&equals_u44;
assign andOp_u61=andOp_u60&port_493b3a04_;
assign equals_u45_a_unsigned=port_77e210a8_;
assign equals_u45_b_unsigned=16'h0;
assign equals_u45=equals_u45_a_unsigned==equals_u45_b_unsigned;
assign lessThan_u25_a_signed=port_1a03f6bd_;
assign lessThan_u25_b_signed=16'h1ff;
assign lessThan_u25=lessThan_u25_a_signed<lessThan_u25_b_signed;
assign andOp_u62=equals_u45&lessThan_u25;
assign equals_u46_a_unsigned=port_1d57b49c_;
assign equals_u46_b_unsigned=32'h20000;
assign equals_u46=equals_u46_a_unsigned==equals_u46_b_unsigned;
assign andOp_u63=andOp_u62&equals_u46;
assign not_u145=!port_493b3a04_;
assign andOp_u64=andOp_u63&not_u145;
assign lessThan_u26_a_unsigned=port_77e210a8_;
assign lessThan_u26_b_unsigned=16'hff;
assign lessThan_u26=lessThan_u26_a_unsigned<lessThan_u26_b_unsigned;
assign lessThan_u27_a_signed=port_1a03f6bd_;
assign lessThan_u27_b_signed=16'h1ff;
assign lessThan_u27=lessThan_u27_a_signed<lessThan_u27_b_signed;
assign andOp_u65=lessThan_u26&lessThan_u27;
assign lessThan_u28_a_unsigned=port_1d57b49c_;
assign lessThan_u28_b_unsigned=32'h20000;
assign lessThan_u28=lessThan_u28_a_unsigned<lessThan_u28_b_unsigned;
assign andOp_u66=andOp_u65&lessThan_u28;
assign andOp_u67=andOp_u66&port_493b3a04_;
assign lessThan_u29_a_unsigned=port_77e210a8_;
assign lessThan_u29_b_unsigned=16'hff;
assign lessThan_u29=lessThan_u29_a_unsigned<lessThan_u29_b_unsigned;
assign lessThan_u30_a_signed=port_1a03f6bd_;
assign lessThan_u30_b_signed=16'h1ff;
assign lessThan_u30=lessThan_u30_a_signed<lessThan_u30_b_signed;
assign andOp_u68=lessThan_u29&lessThan_u30;
assign lessThan_u31_a_unsigned=port_1d57b49c_;
assign lessThan_u31_b_unsigned=32'h20000;
assign lessThan_u31=lessThan_u31_a_unsigned<lessThan_u31_b_unsigned;
assign andOp_u69=andOp_u68&lessThan_u31;
assign not_u146=!port_493b3a04_;
assign andOp_u70=andOp_u69&not_u146;
assign lessThan_u32_a_unsigned=port_77e210a8_;
assign lessThan_u32_b_unsigned=16'hff;
assign lessThan_u32=lessThan_u32_a_unsigned<lessThan_u32_b_unsigned;
assign equals_u47_a_unsigned=port_1d57b49c_;
assign equals_u47_b_unsigned=32'h20000;
assign equals_u47=equals_u47_a_unsigned==equals_u47_b_unsigned;
assign andOp_u71=lessThan_u32&equals_u47;
assign andOp_u72=andOp_u71&port_493b3a04_;
assign lessThan_u33_a_unsigned=port_77e210a8_;
assign lessThan_u33_b_unsigned=16'hff;
assign lessThan_u33=lessThan_u33_a_unsigned<lessThan_u33_b_unsigned;
assign equals_u48_a_unsigned=port_1d57b49c_;
assign equals_u48_b_unsigned=32'h20000;
assign equals_u48=equals_u48_a_unsigned==equals_u48_b_unsigned;
assign andOp_u73=lessThan_u33&equals_u48;
assign not_u147=!port_493b3a04_;
assign andOp_u74=andOp_u73&not_u147;
assign equals_u49_a_unsigned=port_77e210a8_;
assign equals_u49_b_unsigned=16'hff;
assign equals_u49=equals_u49_a_unsigned==equals_u49_b_unsigned;
assign lessThan_u34_a_unsigned=port_1d57b49c_;
assign lessThan_u34_b_unsigned=32'h20000;
assign lessThan_u34=lessThan_u34_a_unsigned<lessThan_u34_b_unsigned;
assign andOp_u75=equals_u49&lessThan_u34;
assign andOp_u76=andOp_u75&port_493b3a04_;
assign equals_u50_a_unsigned=port_77e210a8_;
assign equals_u50_b_unsigned=16'hff;
assign equals_u50=equals_u50_a_unsigned==equals_u50_b_unsigned;
assign lessThan_u35_a_unsigned=port_1d57b49c_;
assign lessThan_u35_b_unsigned=32'h20000;
assign lessThan_u35=lessThan_u35_a_unsigned<lessThan_u35_b_unsigned;
assign andOp_u77=equals_u50&lessThan_u35;
assign not_u148=!port_493b3a04_;
assign andOp_u78=andOp_u77&not_u148;
assign equals_u51_a_unsigned=port_77e210a8_;
assign equals_u51_b_unsigned=16'hff;
assign equals_u51=equals_u51_a_unsigned==equals_u51_b_unsigned;
assign equals_u52_a_unsigned=port_1d57b49c_;
assign equals_u52_b_unsigned=32'h20000;
assign equals_u52=equals_u52_a_unsigned==equals_u52_b_unsigned;
assign andOp_u79=equals_u51&equals_u52;
assign andOp_u80=andOp_u79&port_493b3a04_;
assign equals_u53_a_unsigned=port_77e210a8_;
assign equals_u53_b_unsigned=16'hff;
assign equals_u53=equals_u53_a_unsigned==equals_u53_b_unsigned;
assign equals_u54_a_unsigned=port_1d57b49c_;
assign equals_u54_b_unsigned=32'h20000;
assign equals_u54=equals_u54_a_unsigned==equals_u54_b_unsigned;
assign andOp_u81=equals_u53&equals_u54;
assign not_u149=!port_493b3a04_;
assign andOp_u82=andOp_u81&not_u149;
assign equals_u55_a_unsigned=port_77e210a8_;
assign equals_u55_b_unsigned=16'h0;
assign equals_u55=equals_u55_a_unsigned==equals_u55_b_unsigned;
assign equals_u56_a_signed=port_1a03f6bd_;
assign equals_u56_b_signed=16'h1ff;
assign equals_u56=equals_u56_a_signed==equals_u56_b_signed;
assign andOp_u83=equals_u55&equals_u56;
assign equals_u57_a_unsigned=port_1d57b49c_;
assign equals_u57_b_unsigned=32'h20000;
assign equals_u57=equals_u57_a_unsigned==equals_u57_b_unsigned;
assign andOp_u84=andOp_u83&equals_u57;
assign andOp_u85=andOp_u84&port_493b3a04_;
assign equals_u58_a_unsigned=port_77e210a8_;
assign equals_u58_b_unsigned=16'h0;
assign equals_u58=equals_u58_a_unsigned==equals_u58_b_unsigned;
assign equals_u59_a_signed=port_1a03f6bd_;
assign equals_u59_b_signed=16'h1ff;
assign equals_u59=equals_u59_a_signed==equals_u59_b_signed;
assign andOp_u86=equals_u58&equals_u59;
assign equals_u60_a_unsigned=port_1d57b49c_;
assign equals_u60_b_unsigned=32'h20000;
assign equals_u60=equals_u60_a_unsigned==equals_u60_b_unsigned;
assign andOp_u87=andOp_u86&equals_u60;
assign not_u150=!port_493b3a04_;
assign andOp_u88=andOp_u87&not_u150;
assign lessThan_u36_a_unsigned=port_77e210a8_;
assign lessThan_u36_b_unsigned=16'hff;
assign lessThan_u36=lessThan_u36_a_unsigned<lessThan_u36_b_unsigned;
assign equals_u61_a_unsigned=port_1d57b49c_;
assign equals_u61_b_unsigned=32'h20000;
assign equals_u61=equals_u61_a_unsigned==equals_u61_b_unsigned;
assign andOp_u89=lessThan_u36&equals_u61;
assign andOp_u90=andOp_u89&port_493b3a04_;
assign lessThan_u37_a_unsigned=port_77e210a8_;
assign lessThan_u37_b_unsigned=16'hff;
assign lessThan_u37=lessThan_u37_a_unsigned<lessThan_u37_b_unsigned;
assign equals_u62_a_unsigned=port_1d57b49c_;
assign equals_u62_b_unsigned=32'h20000;
assign equals_u62=equals_u62_a_unsigned==equals_u62_b_unsigned;
assign andOp_u91=lessThan_u37&equals_u62;
assign not_u151=!port_493b3a04_;
assign andOp_u92=andOp_u91&not_u151;
assign equals_u63_a_unsigned=port_77e210a8_;
assign equals_u63_b_unsigned=16'hff;
assign equals_u63=equals_u63_a_unsigned==equals_u63_b_unsigned;
assign equals_u64_a_unsigned=port_1d57b49c_;
assign equals_u64_b_unsigned=32'h20000;
assign equals_u64=equals_u64_a_unsigned==equals_u64_b_unsigned;
assign andOp_u93=equals_u63&equals_u64;
assign andOp_u94=andOp_u93&port_493b3a04_;
assign equals_u65_a_unsigned=port_77e210a8_;
assign equals_u65_b_unsigned=16'hff;
assign equals_u65=equals_u65_a_unsigned==equals_u65_b_unsigned;
assign equals_u66_a_unsigned=port_1d57b49c_;
assign equals_u66_b_unsigned=32'h20000;
assign equals_u66=equals_u66_a_unsigned==equals_u66_b_unsigned;
assign andOp_u95=equals_u65&equals_u66;
assign not_u152=!port_493b3a04_;
assign andOp_u96=andOp_u95&not_u152;
assign equals_u67_a_signed={29'b0, port_2fdf62fc_};
assign equals_u67_b_signed=32'h0;
assign equals_u67=equals_u67_a_signed==equals_u67_b_signed;
assign and_u718_u0=and_u717_u0&not_u153_u0;
assign not_u153_u0=~equals_u67;
assign and_u719_u0=and_u717_u0&equals_u67;
assign andOp_u97=lessThan&port_361addca_;
assign and_u720_u0=and_u727_u0&andOp_u97;
assign and_u721_u0=and_u727_u0&not_u154_u0;
assign not_u154_u0=~andOp_u97;
assign simplePinWrite=and_u725_u0&{1{and_u725_u0}};
assign not_u155_u0=~equals;
assign and_u722_u0=and_u726_u0&equals;
assign and_u723_u0=and_u726_u0&not_u155_u0;
assign simplePinWrite_u123=and_u724_u0&{1{and_u724_u0}};
assign and_u724_u0=and_u722_u0&and_u726_u0;
assign and_u725_u0=and_u720_u0&and_u727_u0;
assign or_u184_u0=and_u725_u0|and_u724_u0;
assign mux_u44=(and_u725_u0)?3'h0:3'h1;
assign and_u726_u0=and_u721_u0&and_u727_u0;
assign and_u727_u0=and_u719_u0&and_u717_u0;
assign equals_u68_a_signed={29'b0, port_2fdf62fc_};
assign equals_u68_b_signed=32'h1;
assign equals_u68=equals_u68_a_signed==equals_u68_b_signed;
assign not_u156_u0=~equals_u68;
assign and_u728_u0=and_u717_u0&equals_u68;
assign and_u729_u0=and_u717_u0&not_u156_u0;
assign not_u157_u0=~port_361addca_;
assign and_u730_u0=and_u738_u0&port_361addca_;
assign and_u731_u0=and_u738_u0&not_u157_u0;
assign and_u732_u0=and_u737_u0&not_u158_u0;
assign and_u733_u0=and_u737_u0&port_687ecc25_;
assign not_u158_u0=~port_687ecc25_;
assign simplePinWrite_u124=and_u734_u0&{1{and_u734_u0}};
assign and_u734_u0=and_u733_u0&and_u737_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_59eedaaa_u0<=1'h0;
else reg_59eedaaa_u0<=and_u735_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_27b4c651_u0<=1'h0;
else reg_27b4c651_u0<=reg_6cac83a7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u35<=1'h0;
else and_delayed_u35<=and_u734_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4a42b705_u0<=1'h0;
else reg_4a42b705_u0<=and_delayed_result_delayed_u3;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_result_delayed_u3<=1'h0;
else and_delayed_result_delayed_u3<=and_delayed_u35;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6cac83a7_u0<=1'h0;
else reg_6cac83a7_u0<=reg_4a42b705_result_delayed_u0;
end
assign or_u185_u0=reg_27b4c651_u0|reg_59eedaaa_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4a42b705_result_delayed_u0<=1'h0;
else reg_4a42b705_result_delayed_u0<=reg_4a42b705_u0;
end
assign and_u735_u0=and_u732_u0&and_u737_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_094d88c9_u0<=1'h0;
else reg_094d88c9_u0<=and_u736_u0;
end
assign and_u736_u0=and_u731_u0&and_u738_u0;
assign or_u186_u0=or_u185_u0|reg_094d88c9_u0;
assign and_u737_u0=and_u730_u0&and_u738_u0;
assign or_u187_u0=or_u186_u0|and_delayed_u36_u0;
assign and_u738_u0=and_u728_u0&and_u717_u0;
assign and_u739_u0=and_u729_u0&and_u717_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u36_u0<=1'h0;
else and_delayed_u36_u0<=and_u739_u0;
end
assign equals_u69_a_signed={29'b0, port_2fdf62fc_};
assign equals_u69_b_signed=32'h2;
assign equals_u69=equals_u69_a_signed==equals_u69_b_signed;
assign and_u740_u0=and_u717_u0&not_u159_u0;
assign not_u159_u0=~equals_u69;
assign and_u741_u0=and_u717_u0&equals_u69;
assign andOp_u98=lessThan_u19&port_361addca_;
assign and_u742_u0=and_u759_u0&not_u160_u0;
assign and_u743_u0=and_u759_u0&andOp_u98;
assign not_u160_u0=~andOp_u98;
assign and_u744_u0=and_u756_u0&not_u161_u0;
assign and_u745_u0=and_u756_u0&port_687ecc25_;
assign not_u161_u0=~port_687ecc25_;
assign simplePinWrite_u125=and_u747_u0&{1{and_u747_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0b7664d7_u0<=1'h0;
else reg_0b7664d7_u0<=and_u747_u0;
end
assign and_u746_u0=and_u744_u0&and_u756_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3ad7a739_u0<=1'h0;
else reg_3ad7a739_u0<=reg_1bc19411_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1bc19411_u0<=1'h0;
else reg_1bc19411_u0<=reg_1b0e6c79_u0;
end
assign and_u747_u0=and_u745_u0&and_u756_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3ad7a739_result_delayed_u0<=1'h0;
else reg_3ad7a739_result_delayed_u0<=reg_3ad7a739_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1b0e6c79_u0<=1'h0;
else reg_1b0e6c79_u0<=reg_0b7664d7_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u37_u0<=1'h0;
else and_delayed_u37_u0<=and_u746_u0;
end
assign or_u188_u0=and_delayed_u37_u0|reg_3ad7a739_result_delayed_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0b7664d7_result_delayed_u0<=1'h0;
else reg_0b7664d7_result_delayed_u0<=reg_0b7664d7_u0;
end
assign andOp_u99=equals_u40&port_361addca_;
assign not_u162_u0=~andOp_u99;
assign and_u748_u0=and_u757_u0&not_u162_u0;
assign and_u749_u0=and_u757_u0&andOp_u99;
assign and_u750_u0=and_u755_u0&not_u163_u0;
assign not_u163_u0=~port_687ecc25_;
assign and_u751_u0=and_u755_u0&port_687ecc25_;
assign simplePinWrite_u126=and_u752_u0&{1{and_u752_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_25e2a223_u0<=1'h0;
else reg_25e2a223_u0<=reg_7132143c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_25e2a223_result_delayed_u0<=1'h0;
else reg_25e2a223_result_delayed_u0<=reg_25e2a223_u0;
end
assign or_u189_u0=reg_25e2a223_result_delayed_u0|and_delayed_u39_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6cb55ed9_u0<=1'h0;
else reg_6cb55ed9_u0<=and_delayed_u38_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7132143c_u0<=1'h0;
else reg_7132143c_u0<=reg_6cb55ed9_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6cb55ed9_result_delayed_u0<=1'h0;
else reg_6cb55ed9_result_delayed_u0<=reg_6cb55ed9_u0;
end
assign and_u752_u0=and_u751_u0&and_u755_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u38_u0<=1'h0;
else and_delayed_u38_u0<=and_u752_u0;
end
assign and_u753_u0=and_u750_u0&and_u755_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u39_u0<=1'h0;
else and_delayed_u39_u0<=and_u753_u0;
end
assign and_u754_u0=and_u748_u0&and_u757_u0;
assign or_u190_u0=or_u189_u0|and_delayed_u40_u0;
assign and_u755_u0=and_u749_u0&and_u757_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u40_u0<=1'h0;
else and_delayed_u40_u0<=and_u754_u0;
end
assign and_u756_u0=and_u743_u0&and_u759_u0;
assign mux_u45_u0=(and_u747_u0)?3'h2:3'h3;
assign or_u191_u0=and_u747_u0|and_u752_u0;
assign or_u192_u0=or_u190_u0|or_u188_u0;
assign and_u757_u0=and_u742_u0&and_u759_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_43562f66_u0<=1'h0;
else reg_43562f66_u0<=and_u758_u0;
end
assign or_u193_u0=or_u192_u0|reg_43562f66_u0;
assign and_u758_u0=and_u740_u0&and_u717_u0;
assign and_u759_u0=and_u741_u0&and_u717_u0;
assign equals_u70_a_signed={29'b0, port_2fdf62fc_};
assign equals_u70_b_signed=32'h3;
assign equals_u70=equals_u70_a_signed==equals_u70_b_signed;
assign not_u164_u0=~equals_u70;
assign and_u760_u0=and_u717_u0&not_u164_u0;
assign and_u761_u0=and_u717_u0&equals_u70;
assign andOp_u100=andOp_u55&port_361addca_;
assign not_u165_u0=~andOp_u100;
assign and_u762_u0=and_u794_u0&andOp_u100;
assign and_u763_u0=and_u794_u0&not_u165_u0;
assign and_u764_u0=and_u793_u0&port_687ecc25_;
assign and_u765_u0=and_u793_u0&not_u166_u0;
assign not_u166_u0=~port_687ecc25_;
assign simplePinWrite_u127=and_u767_u0&{1{and_u767_u0}};
assign and_u766_u0=and_u765_u0&and_u793_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6f936df5_u0<=1'h0;
else reg_6f936df5_u0<=reg_5373c17a_result_delayed_u0;
end
assign or_u194_u0=reg_6f936df5_result_delayed_result_delayed_result_delayed_u0|and_delayed_u41_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5373c17a_u0<=1'h0;
else reg_5373c17a_u0<=and_u767_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5373c17a_result_delayed_u0<=1'h0;
else reg_5373c17a_result_delayed_u0<=reg_5373c17a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u41_u0<=1'h0;
else and_delayed_u41_u0<=and_u766_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6f936df5_result_delayed_u0<=1'h0;
else reg_6f936df5_result_delayed_u0<=reg_6f936df5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6f936df5_result_delayed_result_delayed_u0<=1'h0;
else reg_6f936df5_result_delayed_result_delayed_u0<=reg_6f936df5_result_delayed_u0;
end
assign and_u767_u0=and_u764_u0&and_u793_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6f936df5_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_6f936df5_result_delayed_result_delayed_result_delayed_u0<=reg_6f936df5_result_delayed_result_delayed_u0;
end
assign andOp_u101=andOp_u58&port_361addca_;
assign and_u768_u0=and_u792_u0&not_u167_u0;
assign not_u167_u0=~andOp_u101;
assign and_u769_u0=and_u792_u0&andOp_u101;
assign and_u770_u0=and_u790_u0&port_4533a20c_;
assign not_u168_u0=~port_4533a20c_;
assign and_u771_u0=and_u790_u0&not_u168_u0;
assign simplePinWrite_u128=and_u772_u0&{1{and_u772_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_74073fe4_u0<=1'h0;
else reg_74073fe4_u0<=and_u773_u0;
end
assign and_u772_u0=and_u770_u0&and_u790_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0eaacf63_u0<=1'h0;
else reg_0eaacf63_u0<=reg_3acc3e9c_u0;
end
assign or_u195_u0=reg_74073fe4_u0|reg_24425050_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u42_u0<=1'h0;
else and_delayed_u42_u0<=and_u772_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3acc3e9c_u0<=1'h0;
else reg_3acc3e9c_u0<=and_delayed_result_delayed_u4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_24425050_u0<=1'h0;
else reg_24425050_u0<=reg_0eaacf63_result_delayed_u0;
end
assign and_u773_u0=and_u771_u0&and_u790_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_result_delayed_u4_u0<=1'h0;
else and_delayed_result_delayed_u4_u0<=and_delayed_u42_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0eaacf63_result_delayed_u0<=1'h0;
else reg_0eaacf63_result_delayed_u0<=reg_0eaacf63_u0;
end
assign and_u774_u0=and_u791_u0&andOp_u61;
assign and_u775_u0=and_u791_u0&not_u169_u0;
assign not_u169_u0=~andOp_u61;
assign and_u776_u0=and_u789_u0&port_687ecc25_;
assign and_u777_u0=and_u789_u0&not_u170_u0;
assign not_u170_u0=~port_687ecc25_;
assign simplePinWrite_u129=and_u778_u0&{1{and_u778_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_774e2f4e_u0<=1'h0;
else reg_774e2f4e_u0<=reg_376a948f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1efbe559_u0<=1'h0;
else reg_1efbe559_u0<=and_u779_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_376a948f_u0<=1'h0;
else reg_376a948f_u0<=and_delayed_u43_u0;
end
assign and_u778_u0=and_u776_u0&and_u789_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4094683f_u0<=1'h0;
else reg_4094683f_u0<=reg_774e2f4e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_774e2f4e_result_delayed_u0<=1'h0;
else reg_774e2f4e_result_delayed_u0<=reg_774e2f4e_u0;
end
assign or_u196_u0=reg_4094683f_u0|reg_1efbe559_u0;
assign and_u779_u0=and_u777_u0&and_u789_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u43_u0<=1'h0;
else and_delayed_u43_u0<=and_u778_u0;
end
assign and_u780_u0=and_u788_u0&not_u171_u0;
assign and_u781_u0=and_u788_u0&andOp_u64;
assign not_u171_u0=~andOp_u64;
assign and_u782_u0=and_u787_u0&port_4533a20c_;
assign and_u783_u0=and_u787_u0&not_u172_u0;
assign not_u172_u0=~port_4533a20c_;
assign simplePinWrite_u130=and_u785_u0&{1{and_u785_u0}};
assign and_u784_u0=and_u783_u0&and_u787_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_549c7b3d_u0<=1'h0;
else reg_549c7b3d_u0<=and_u785_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3da7ac05_u0<=1'h0;
else reg_3da7ac05_u0<=reg_549c7b3d_result_delayed_u0;
end
assign or_u197_u0=and_delayed_u44_u0|reg_3da7ac05_result_delayed_result_delayed_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u44_u0<=1'h0;
else and_delayed_u44_u0<=and_u784_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_549c7b3d_result_delayed_u0<=1'h0;
else reg_549c7b3d_result_delayed_u0<=reg_549c7b3d_u0;
end
assign and_u785_u0=and_u782_u0&and_u787_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3da7ac05_result_delayed_u0<=1'h0;
else reg_3da7ac05_result_delayed_u0<=reg_3da7ac05_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3da7ac05_result_delayed_result_delayed_u0<=1'h0;
else reg_3da7ac05_result_delayed_result_delayed_u0<=reg_3da7ac05_result_delayed_u0;
end
assign and_u786_u0=and_u780_u0&and_u788_u0;
assign or_u198_u0=or_u197_u0|and_delayed_u45_u0;
assign and_u787_u0=and_u781_u0&and_u788_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u45_u0<=1'h0;
else and_delayed_u45_u0<=and_u786_u0;
end
assign or_u199_u0=or_u196_u0|or_u198_u0;
assign or_u200_u0=and_u778_u0|and_u785_u0;
assign and_u788_u0=and_u775_u0&and_u791_u0;
assign and_u789_u0=and_u774_u0&and_u791_u0;
assign or_u201_u0=and_u772_u0|or_u200_u0;
assign and_u790_u0=and_u769_u0&and_u792_u0;
assign or_u202_u0=or_u199_u0|or_u195_u0;
assign and_u791_u0=and_u768_u0&and_u792_u0;
assign or_u203_u0=or_u194_u0|or_u202_u0;
assign or_u204_u0=and_u767_u0|or_u201_u0;
assign and_u792_u0=and_u763_u0&and_u794_u0;
assign and_u793_u0=and_u762_u0&and_u794_u0;
assign or_u205_u0=or_u203_u0|reg_05c7e893_u0;
assign and_u794_u0=and_u761_u0&and_u717_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_05c7e893_u0<=1'h0;
else reg_05c7e893_u0<=and_u795_u0;
end
assign and_u795_u0=and_u760_u0&and_u717_u0;
assign equals_u71_a_signed={29'b0, port_2fdf62fc_};
assign equals_u71_b_signed=32'h4;
assign equals_u71=equals_u71_a_signed==equals_u71_b_signed;
assign and_u796_u0=and_u717_u0&not_u173_u0;
assign not_u173_u0=~equals_u71;
assign and_u797_u0=and_u717_u0&equals_u71;
assign andOp_u102=andOp_u67&port_361addca_;
assign and_u798_u0=and_u862_u0&not_u174_u0;
assign and_u799_u0=and_u862_u0&andOp_u102;
assign not_u174_u0=~andOp_u102;
assign and_u800_u0=and_u860_u0&port_687ecc25_;
assign and_u801_u0=and_u860_u0&not_u175_u0;
assign not_u175_u0=~port_687ecc25_;
assign simplePinWrite_u131=and_u803_u0&{1{and_u803_u0}};
assign or_u206_u0=reg_74ec09a7_u0|and_delayed_u46_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3226eb2c_u0<=1'h0;
else reg_3226eb2c_u0<=and_u803_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_23c4568f_u0<=1'h0;
else reg_23c4568f_u0<=reg_648fa1fc_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_74ec09a7_u0<=1'h0;
else reg_74ec09a7_u0<=reg_23c4568f_result_delayed_u0;
end
assign and_u802_u0=and_u801_u0&and_u860_u0;
assign and_u803_u0=and_u800_u0&and_u860_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_23c4568f_result_delayed_u0<=1'h0;
else reg_23c4568f_result_delayed_u0<=reg_23c4568f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_648fa1fc_u0<=1'h0;
else reg_648fa1fc_u0<=reg_3226eb2c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u46_u0<=1'h0;
else and_delayed_u46_u0<=and_u802_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3226eb2c_result_delayed_u0<=1'h0;
else reg_3226eb2c_result_delayed_u0<=reg_3226eb2c_u0;
end
assign andOp_u103=andOp_u70&port_361addca_;
assign not_u176_u0=~andOp_u103;
assign and_u804_u0=and_u861_u0&andOp_u103;
assign and_u805_u0=and_u861_u0&not_u176_u0;
assign and_u806_u0=and_u858_u0&port_4533a20c_;
assign not_u177_u0=~port_4533a20c_;
assign and_u807_u0=and_u858_u0&not_u177_u0;
assign simplePinWrite_u132=and_u808_u0&{1{and_u808_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4fea946b_u0<=1'h0;
else reg_4fea946b_u0<=and_delayed_u47_u0;
end
assign and_u808_u0=and_u806_u0&and_u858_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6e00556b_u0<=1'h0;
else reg_6e00556b_u0<=reg_309dfcec_u0;
end
assign or_u207_u0=reg_7b04c971_u0|reg_6e00556b_result_delayed_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6e00556b_result_delayed_u0<=1'h0;
else reg_6e00556b_result_delayed_u0<=reg_6e00556b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_309dfcec_u0<=1'h0;
else reg_309dfcec_u0<=reg_4fea946b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u47_u0<=1'h0;
else and_delayed_u47_u0<=and_u808_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7b04c971_u0<=1'h0;
else reg_7b04c971_u0<=and_u809_u0;
end
assign and_u809_u0=and_u807_u0&and_u858_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4fea946b_result_delayed_u0<=1'h0;
else reg_4fea946b_result_delayed_u0<=reg_4fea946b_u0;
end
assign not_u178_u0=~andOp_u72;
assign and_u810_u0=and_u859_u0&andOp_u72;
assign and_u811_u0=and_u859_u0&not_u178_u0;
assign not_u179_u0=~port_687ecc25_;
assign and_u812_u0=and_u856_u0&not_u179_u0;
assign and_u813_u0=and_u856_u0&port_687ecc25_;
assign simplePinWrite_u133=and_u815_u0&{1{and_u815_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7cdd073f_u0<=1'h0;
else reg_7cdd073f_u0<=and_u815_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01b946ba_u0<=1'h0;
else reg_01b946ba_u0<=reg_526cf179_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01b946ba_result_delayed_u0<=1'h0;
else reg_01b946ba_result_delayed_u0<=reg_01b946ba_u0;
end
assign and_u814_u0=and_u812_u0&and_u856_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_526cf179_u0<=1'h0;
else reg_526cf179_u0<=reg_7cdd073f_result_delayed_u0;
end
assign or_u208_u0=reg_01b946ba_result_delayed_u0|and_delayed_u48_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u48_u0<=1'h0;
else and_delayed_u48_u0<=and_u814_u0;
end
assign and_u815_u0=and_u813_u0&and_u856_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7cdd073f_result_delayed_u0<=1'h0;
else reg_7cdd073f_result_delayed_u0<=reg_7cdd073f_u0;
end
assign and_u816_u0=and_u857_u0&andOp_u74;
assign not_u180_u0=~andOp_u74;
assign and_u817_u0=and_u857_u0&not_u180_u0;
assign and_u818_u0=and_u854_u0&port_4533a20c_;
assign and_u819_u0=and_u854_u0&not_u181_u0;
assign not_u181_u0=~port_4533a20c_;
assign simplePinWrite_u134=and_u821_u0&{1{and_u821_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_49ca584b_u0<=1'h0;
else reg_49ca584b_u0<=reg_033b743f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_033b743f_u0<=1'h0;
else reg_033b743f_u0<=and_delayed_u50_u0;
end
assign and_u820_u0=and_u819_u0&and_u854_u0;
assign or_u209_u0=and_delayed_u49_u0|reg_49ca584b_result_delayed_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u49_u0<=1'h0;
else and_delayed_u49_u0<=and_u820_u0;
end
assign and_u821_u0=and_u818_u0&and_u854_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_033b743f_result_delayed_u0<=1'h0;
else reg_033b743f_result_delayed_u0<=reg_033b743f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u50_u0<=1'h0;
else and_delayed_u50_u0<=and_u821_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_49ca584b_result_delayed_u0<=1'h0;
else reg_49ca584b_result_delayed_u0<=reg_49ca584b_u0;
end
assign andOp_u104=andOp_u76&port_361addca_;
assign and_u822_u0=and_u855_u0&andOp_u104;
assign and_u823_u0=and_u855_u0&not_u182_u0;
assign not_u182_u0=~andOp_u104;
assign not_u183_u0=~port_687ecc25_;
assign and_u824_u0=and_u853_u0&port_687ecc25_;
assign and_u825_u0=and_u853_u0&not_u183_u0;
assign simplePinWrite_u135=and_u827_u0&{1{and_u827_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_38c345e9_u0<=1'h0;
else reg_38c345e9_u0<=and_u827_u0;
end
assign and_u826_u0=and_u825_u0&and_u853_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0d74457a_u0<=1'h0;
else reg_0d74457a_u0<=reg_2f356d21_u0;
end
assign and_u827_u0=and_u824_u0&and_u853_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2f356d21_u0<=1'h0;
else reg_2f356d21_u0<=reg_38c345e9_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u51_u0<=1'h0;
else and_delayed_u51_u0<=and_u826_u0;
end
assign or_u210_u0=and_delayed_u51_u0|reg_0d74457a_result_delayed_result_delayed_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_38c345e9_result_delayed_u0<=1'h0;
else reg_38c345e9_result_delayed_u0<=reg_38c345e9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0d74457a_result_delayed_u0<=1'h0;
else reg_0d74457a_result_delayed_u0<=reg_0d74457a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0d74457a_result_delayed_result_delayed_u0<=1'h0;
else reg_0d74457a_result_delayed_result_delayed_u0<=reg_0d74457a_result_delayed_u0;
end
assign andOp_u105=andOp_u78&port_361addca_;
assign not_u184_u0=~andOp_u105;
assign and_u828_u0=and_u852_u0&andOp_u105;
assign and_u829_u0=and_u852_u0&not_u184_u0;
assign not_u185_u0=~port_4533a20c_;
assign and_u830_u0=and_u851_u0&port_4533a20c_;
assign and_u831_u0=and_u851_u0&not_u185_u0;
assign simplePinWrite_u136=and_u833_u0&{1{and_u833_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_317cd17d_u0<=1'h0;
else reg_317cd17d_u0<=and_delayed_u52_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_002dc3a9_u0<=1'h0;
else reg_002dc3a9_u0<=and_u832_u0;
end
assign or_u211_u0=reg_002dc3a9_u0|reg_624de640_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_71ed30e6_u0<=1'h0;
else reg_71ed30e6_u0<=reg_317cd17d_result_delayed_u0;
end
assign and_u832_u0=and_u831_u0&and_u851_u0;
assign and_u833_u0=and_u830_u0&and_u851_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_624de640_u0<=1'h0;
else reg_624de640_u0<=reg_71ed30e6_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_317cd17d_result_delayed_u0<=1'h0;
else reg_317cd17d_result_delayed_u0<=reg_317cd17d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u52_u0<=1'h0;
else and_delayed_u52_u0<=and_u833_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_71ed30e6_result_delayed_u0<=1'h0;
else reg_71ed30e6_result_delayed_u0<=reg_71ed30e6_u0;
end
assign and_u834_u0=and_u850_u0&andOp_u80;
assign not_u186_u0=~andOp_u80;
assign and_u835_u0=and_u850_u0&not_u186_u0;
assign and_u836_u0=and_u849_u0&not_u187_u0;
assign not_u187_u0=~port_687ecc25_;
assign and_u837_u0=and_u849_u0&port_687ecc25_;
assign simplePinWrite_u137=and_u838_u0&{1{and_u838_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_63fb95d2_u0<=1'h0;
else reg_63fb95d2_u0<=reg_398c8621_u0;
end
assign or_u212_u0=reg_63fb95d2_result_delayed_result_delayed_u0|reg_4529a71b_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_398c8621_u0<=1'h0;
else reg_398c8621_u0<=and_delayed_u53_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_63fb95d2_result_delayed_u0<=1'h0;
else reg_63fb95d2_result_delayed_u0<=reg_63fb95d2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_63fb95d2_result_delayed_result_delayed_u0<=1'h0;
else reg_63fb95d2_result_delayed_result_delayed_u0<=reg_63fb95d2_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4529a71b_u0<=1'h0;
else reg_4529a71b_u0<=and_u839_u0;
end
assign and_u838_u0=and_u837_u0&and_u849_u0;
assign and_u839_u0=and_u836_u0&and_u849_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u53_u0<=1'h0;
else and_delayed_u53_u0<=and_u838_u0;
end
assign and_u840_u0=and_u848_u0&not_u188_u0;
assign and_u841_u0=and_u848_u0&andOp_u82;
assign not_u188_u0=~andOp_u82;
assign and_u842_u0=and_u847_u0&not_u189_u0;
assign and_u843_u0=and_u847_u0&port_4533a20c_;
assign not_u189_u0=~port_4533a20c_;
assign simplePinWrite_u138=and_u844_u0&{1{and_u844_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_420f216e_u0<=1'h0;
else reg_420f216e_u0<=reg_6e40f982_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6e40f982_u0<=1'h0;
else reg_6e40f982_u0<=reg_15a02ae4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2d931bb0_u0<=1'h0;
else reg_2d931bb0_u0<=and_u844_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_15a02ae4_u0<=1'h0;
else reg_15a02ae4_u0<=reg_2d931bb0_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3b71b3f6_u0<=1'h0;
else reg_3b71b3f6_u0<=and_u845_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2d931bb0_result_delayed_u0<=1'h0;
else reg_2d931bb0_result_delayed_u0<=reg_2d931bb0_u0;
end
assign or_u213_u0=reg_420f216e_u0|reg_3b71b3f6_u0;
assign and_u844_u0=and_u843_u0&and_u847_u0;
assign and_u845_u0=and_u842_u0&and_u847_u0;
assign and_u846_u0=and_u840_u0&and_u848_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u54_u0<=1'h0;
else and_delayed_u54_u0<=and_u846_u0;
end
assign and_u847_u0=and_u841_u0&and_u848_u0;
assign or_u214_u0=and_delayed_u54_u0|or_u213_u0;
assign or_u215_u0=or_u212_u0|or_u214_u0;
assign or_u216_u0=and_u838_u0|and_u844_u0;
assign and_u848_u0=and_u835_u0&and_u850_u0;
assign and_u849_u0=and_u834_u0&and_u850_u0;
assign or_u217_u0=or_u215_u0|or_u211_u0;
assign or_u218_u0=and_u833_u0|or_u216_u0;
assign and_u850_u0=and_u829_u0&and_u852_u0;
assign and_u851_u0=and_u828_u0&and_u852_u0;
assign and_u852_u0=and_u823_u0&and_u855_u0;
assign or_u219_u0=or_u210_u0|or_u217_u0;
assign or_u220_u0=and_u827_u0|or_u218_u0;
assign and_u853_u0=and_u822_u0&and_u855_u0;
assign and_u854_u0=and_u816_u0&and_u857_u0;
assign or_u221_u0=or_u209_u0|or_u219_u0;
assign mux_u46_u0=(and_u821_u0)?3'h4:3'h5;
assign or_u222_u0=and_u821_u0|or_u220_u0;
assign and_u855_u0=and_u817_u0&and_u857_u0;
assign or_u223_u0=or_u208_u0|or_u221_u0;
assign and_u856_u0=and_u810_u0&and_u859_u0;
assign and_u857_u0=and_u811_u0&and_u859_u0;
assign mux_u47_u0=(and_u815_u0)?3'h4:{2'b10, mux_u46_u0[0]};
assign or_u224_u0=and_u815_u0|or_u222_u0;
assign and_u858_u0=and_u804_u0&and_u861_u0;
assign or_u225_u0=or_u223_u0|or_u207_u0;
assign or_u226_u0=and_u808_u0|or_u224_u0;
assign mux_u48_u0=(and_u808_u0)?3'h4:{2'b10, mux_u47_u0[0]};
assign and_u859_u0=and_u805_u0&and_u861_u0;
assign mux_u49_u0=(and_u803_u0)?3'h4:{2'b10, mux_u48_u0[0]};
assign or_u227_u0=and_u803_u0|or_u226_u0;
assign and_u860_u0=and_u799_u0&and_u862_u0;
assign or_u228_u0=or_u225_u0|or_u206_u0;
assign and_u861_u0=and_u798_u0&and_u862_u0;
assign and_u862_u0=and_u797_u0&and_u717_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_17b91f93_u0<=1'h0;
else reg_17b91f93_u0<=and_u863_u0;
end
assign or_u229_u0=or_u228_u0|reg_17b91f93_u0;
assign and_u863_u0=and_u796_u0&and_u717_u0;
assign equals_u72_a_signed={29'b0, port_2fdf62fc_};
assign equals_u72_b_signed=32'h5;
assign equals_u72=equals_u72_a_signed==equals_u72_b_signed;
assign and_u864_u0=and_u717_u0&equals_u72;
assign not_u190_u0=~equals_u72;
assign and_u865_u0=and_u717_u0&not_u190_u0;
assign andOp_u106=andOp_u55&port_361addca_;
assign and_u866_u0=and_u915_u0&not_u191_u0;
assign and_u867_u0=and_u915_u0&andOp_u106;
assign not_u191_u0=~andOp_u106;
assign not_u192_u0=~port_687ecc25_;
assign and_u868_u0=and_u912_u0&port_687ecc25_;
assign and_u869_u0=and_u912_u0&not_u192_u0;
assign simplePinWrite_u139=and_u871_u0&{1{and_u871_u0}};
assign and_u870_u0=and_u869_u0&and_u912_u0;
assign and_u871_u0=and_u868_u0&and_u912_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_62867c89_u0<=1'h0;
else reg_62867c89_u0<=reg_342b0dff_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u55_u0<=1'h0;
else and_delayed_u55_u0<=and_u871_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_342b0dff_u0<=1'h0;
else reg_342b0dff_u0<=and_delayed_result_delayed_u5_u0;
end
assign or_u230_u0=reg_62867c89_result_delayed_u0|and_delayed_u56_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_342b0dff_result_delayed_u0<=1'h0;
else reg_342b0dff_result_delayed_u0<=reg_342b0dff_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_62867c89_result_delayed_u0<=1'h0;
else reg_62867c89_result_delayed_u0<=reg_62867c89_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_result_delayed_u5_u0<=1'h0;
else and_delayed_result_delayed_u5_u0<=and_delayed_u55_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u56_u0<=1'h0;
else and_delayed_u56_u0<=and_u870_u0;
end
assign andOp_u107=andOp_u58&port_361addca_;
assign not_u193_u0=~andOp_u107;
assign and_u872_u0=and_u913_u0&andOp_u107;
assign and_u873_u0=and_u913_u0&not_u193_u0;
assign and_u874_u0=and_u911_u0&port_4533a20c_;
assign and_u875_u0=and_u911_u0&not_u194_u0;
assign not_u194_u0=~port_4533a20c_;
assign simplePinWrite_u140=and_u877_u0&{1{and_u877_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5c254b63_u0<=1'h0;
else reg_5c254b63_u0<=reg_4dcbcd47_result_delayed_u0;
end
assign and_u876_u0=and_u875_u0&and_u911_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_122ac30d_u0<=1'h0;
else reg_122ac30d_u0<=reg_5c254b63_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4dcbcd47_u0<=1'h0;
else reg_4dcbcd47_u0<=and_delayed_u58_u0;
end
assign and_u877_u0=and_u874_u0&and_u911_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5c254b63_result_delayed_u0<=1'h0;
else reg_5c254b63_result_delayed_u0<=reg_5c254b63_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u57_u0<=1'h0;
else and_delayed_u57_u0<=and_u876_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4dcbcd47_result_delayed_u0<=1'h0;
else reg_4dcbcd47_result_delayed_u0<=reg_4dcbcd47_u0;
end
assign or_u231_u0=reg_122ac30d_u0|and_delayed_u57_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u58_u0<=1'h0;
else and_delayed_u58_u0<=and_u877_u0;
end
assign not_u195_u0=~andOp_u61;
assign and_u878_u0=and_u910_u0&andOp_u61;
assign and_u879_u0=and_u910_u0&not_u195_u0;
assign and_u880_u0=and_u909_u0&port_687ecc25_;
assign and_u881_u0=and_u909_u0&not_u196_u0;
assign not_u196_u0=~port_687ecc25_;
assign simplePinWrite_u141=and_u883_u0&{1{and_u883_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4aef9f0e_u0<=1'h0;
else reg_4aef9f0e_u0<=reg_307315fd_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_77e48187_u0<=1'h0;
else reg_77e48187_u0<=and_u882_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4aef9f0e_result_delayed_u0<=1'h0;
else reg_4aef9f0e_result_delayed_u0<=reg_4aef9f0e_u0;
end
assign or_u232_u0=reg_77e48187_u0|reg_4aef9f0e_result_delayed_result_delayed_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_307315fd_u0<=1'h0;
else reg_307315fd_u0<=and_u883_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_307315fd_result_delayed_u0<=1'h0;
else reg_307315fd_result_delayed_u0<=reg_307315fd_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4aef9f0e_result_delayed_result_delayed_u0<=1'h0;
else reg_4aef9f0e_result_delayed_result_delayed_u0<=reg_4aef9f0e_result_delayed_u0;
end
assign and_u882_u0=and_u881_u0&and_u909_u0;
assign and_u883_u0=and_u880_u0&and_u909_u0;
assign and_u884_u0=and_u908_u0&not_u197_u0;
assign not_u197_u0=~andOp_u64;
assign and_u885_u0=and_u908_u0&andOp_u64;
assign and_u886_u0=and_u906_u0&not_u198_u0;
assign and_u887_u0=and_u906_u0&port_4533a20c_;
assign not_u198_u0=~port_4533a20c_;
assign simplePinWrite_u142=and_u888_u0&{1{and_u888_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7ee43ce2_u0<=1'h0;
else reg_7ee43ce2_u0<=and_delayed_u59_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_32619689_u0<=1'h0;
else reg_32619689_u0<=reg_7ee43ce2_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5416fdbe_u0<=1'h0;
else reg_5416fdbe_u0<=and_u889_u0;
end
assign or_u233_u0=reg_32619689_result_delayed_u0|reg_5416fdbe_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_32619689_result_delayed_u0<=1'h0;
else reg_32619689_result_delayed_u0<=reg_32619689_u0;
end
assign and_u888_u0=and_u887_u0&and_u906_u0;
assign and_u889_u0=and_u886_u0&and_u906_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7ee43ce2_result_delayed_u0<=1'h0;
else reg_7ee43ce2_result_delayed_u0<=reg_7ee43ce2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u59_u0<=1'h0;
else and_delayed_u59_u0<=and_u888_u0;
end
assign not_u199_u0=~andOp_u85;
assign and_u890_u0=and_u907_u0&andOp_u85;
assign and_u891_u0=and_u907_u0&not_u199_u0;
assign and_u892_u0=and_u905_u0&port_687ecc25_;
assign and_u893_u0=and_u905_u0&not_u200_u0;
assign not_u200_u0=~port_687ecc25_;
assign simplePinWrite_u143=and_u894_u0&{1{and_u894_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a4edfae_u0<=1'h0;
else reg_7a4edfae_u0<=reg_25cc270d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_25cc270d_u0<=1'h0;
else reg_25cc270d_u0<=reg_5b6f804b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5b6f804b_u0<=1'h0;
else reg_5b6f804b_u0<=and_delayed_result_delayed_u6_u0;
end
assign and_u894_u0=and_u892_u0&and_u905_u0;
assign and_u895_u0=and_u893_u0&and_u905_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u60_u0<=1'h0;
else and_delayed_u60_u0<=and_u894_u0;
end
assign or_u234_u0=reg_7a4edfae_u0|and_delayed_u61_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u61_u0<=1'h0;
else and_delayed_u61_u0<=and_u895_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_result_delayed_u6_u0<=1'h0;
else and_delayed_result_delayed_u6_u0<=and_delayed_u60_u0;
end
assign and_u896_u0=and_u904_u0&not_u201_u0;
assign not_u201_u0=~andOp_u88;
assign and_u897_u0=and_u904_u0&andOp_u88;
assign and_u898_u0=and_u902_u0&not_u202_u0;
assign not_u202_u0=~port_4533a20c_;
assign and_u899_u0=and_u902_u0&port_4533a20c_;
assign simplePinWrite_u144=and_u901_u0&{1{and_u901_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_07a24aa2_u0<=1'h0;
else reg_07a24aa2_u0<=reg_5887a60e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5887a60e_u0<=1'h0;
else reg_5887a60e_u0<=and_u901_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0281fc6b_u0<=1'h0;
else reg_0281fc6b_u0<=reg_07a24aa2_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0281fc6b_result_delayed_u0<=1'h0;
else reg_0281fc6b_result_delayed_u0<=reg_0281fc6b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_07a24aa2_result_delayed_u0<=1'h0;
else reg_07a24aa2_result_delayed_u0<=reg_07a24aa2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_09dc81cd_u0<=1'h0;
else reg_09dc81cd_u0<=and_u900_u0;
end
assign and_u900_u0=and_u898_u0&and_u902_u0;
assign and_u901_u0=and_u899_u0&and_u902_u0;
assign or_u235_u0=reg_0281fc6b_result_delayed_u0|reg_09dc81cd_u0;
assign and_u902_u0=and_u897_u0&and_u904_u0;
assign and_u903_u0=and_u896_u0&and_u904_u0;
assign or_u236_u0=or_u235_u0|and_delayed_u62_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u62_u0<=1'h0;
else and_delayed_u62_u0<=and_u903_u0;
end
assign and_u904_u0=and_u891_u0&and_u907_u0;
assign or_u237_u0=and_u894_u0|and_u901_u0;
assign and_u905_u0=and_u890_u0&and_u907_u0;
assign or_u238_u0=or_u236_u0|or_u234_u0;
assign and_u906_u0=and_u885_u0&and_u908_u0;
assign mux_u50_u0=(and_u888_u0)?3'h4:3'h6;
assign or_u239_u0=and_u888_u0|or_u237_u0;
assign and_u907_u0=and_u884_u0&and_u908_u0;
assign or_u240_u0=or_u233_u0|or_u238_u0;
assign and_u908_u0=and_u879_u0&and_u910_u0;
assign or_u241_u0=or_u232_u0|or_u240_u0;
assign and_u909_u0=and_u878_u0&and_u910_u0;
assign mux_u51_u0=(and_u883_u0)?3'h4:{1'b1, mux_u50_u0[1], 1'b0};
assign or_u242_u0=and_u883_u0|or_u239_u0;
assign and_u910_u0=and_u873_u0&and_u913_u0;
assign and_u911_u0=and_u872_u0&and_u913_u0;
assign or_u243_u0=or_u231_u0|or_u241_u0;
assign mux_u52_u0=(and_u877_u0)?3'h4:{1'b1, mux_u51_u0[1], 1'b0};
assign or_u244_u0=and_u877_u0|or_u242_u0;
assign and_u912_u0=and_u867_u0&and_u915_u0;
assign or_u245_u0=or_u243_u0|or_u230_u0;
assign mux_u53_u0=(and_u871_u0)?3'h4:{1'b1, mux_u52_u0[1], 1'b0};
assign or_u246_u0=and_u871_u0|or_u244_u0;
assign and_u913_u0=and_u866_u0&and_u915_u0;
assign or_u247_u0=or_u245_u0|and_delayed_u63_u0;
assign and_u914_u0=and_u865_u0&and_u717_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u63_u0<=1'h0;
else and_delayed_u63_u0<=and_u914_u0;
end
assign and_u915_u0=and_u864_u0&and_u717_u0;
assign equals_u73_a_signed={29'b0, port_2fdf62fc_};
assign equals_u73_b_signed=32'h6;
assign equals_u73=equals_u73_a_signed==equals_u73_b_signed;
assign and_u916_u0=and_u717_u0&equals_u73;
assign not_u203_u0=~equals_u73;
assign and_u917_u0=and_u717_u0&not_u203_u0;
assign and_u918_u0=and_u950_u0&not_u204_u0;
assign not_u204_u0=~andOp_u90;
assign and_u919_u0=and_u950_u0&andOp_u90;
assign and_u920_u0=and_u949_u0&port_687ecc25_;
assign not_u205_u0=~port_687ecc25_;
assign and_u921_u0=and_u949_u0&not_u205_u0;
assign simplePinWrite_u145=and_u923_u0&{1{and_u923_u0}};
assign and_u922_u0=and_u921_u0&and_u949_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5938427c_u0<=1'h0;
else reg_5938427c_u0<=reg_3a61ec86_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3a61ec86_u0<=1'h0;
else reg_3a61ec86_u0<=and_delayed_u65_u0;
end
assign and_u923_u0=and_u920_u0&and_u949_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u64_u0<=1'h0;
else and_delayed_u64_u0<=and_u922_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u65_u0<=1'h0;
else and_delayed_u65_u0<=and_u923_u0;
end
assign or_u248_u0=reg_5938427c_result_delayed_result_delayed_u0|and_delayed_u64_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5938427c_result_delayed_u0<=1'h0;
else reg_5938427c_result_delayed_u0<=reg_5938427c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5938427c_result_delayed_result_delayed_u0<=1'h0;
else reg_5938427c_result_delayed_result_delayed_u0<=reg_5938427c_result_delayed_u0;
end
assign and_u924_u0=and_u948_u0&not_u206_u0;
assign and_u925_u0=and_u948_u0&andOp_u92;
assign not_u206_u0=~andOp_u92;
assign not_u207_u0=~port_4533a20c_;
assign and_u926_u0=and_u947_u0&port_4533a20c_;
assign and_u927_u0=and_u947_u0&not_u207_u0;
assign simplePinWrite_u146=and_u928_u0&{1{and_u928_u0}};
assign and_u928_u0=and_u926_u0&and_u947_u0;
assign or_u249_u0=reg_5a1c7caf_u0|reg_0c3b0433_result_delayed_result_delayed_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0c3b0433_u0<=1'h0;
else reg_0c3b0433_u0<=and_delayed_result_delayed_u7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u66_u0<=1'h0;
else and_delayed_u66_u0<=and_u928_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5a1c7caf_u0<=1'h0;
else reg_5a1c7caf_u0<=and_u929_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_result_delayed_u7_u0<=1'h0;
else and_delayed_result_delayed_u7_u0<=and_delayed_u66_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0c3b0433_result_delayed_u0<=1'h0;
else reg_0c3b0433_result_delayed_u0<=reg_0c3b0433_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0c3b0433_result_delayed_result_delayed_u0<=1'h0;
else reg_0c3b0433_result_delayed_result_delayed_u0<=reg_0c3b0433_result_delayed_u0;
end
assign and_u929_u0=and_u927_u0&and_u947_u0;
assign not_u208_u0=~andOp_u94;
assign and_u930_u0=and_u946_u0&andOp_u94;
assign and_u931_u0=and_u946_u0&not_u208_u0;
assign and_u932_u0=and_u945_u0&port_687ecc25_;
assign and_u933_u0=and_u945_u0&not_u209_u0;
assign not_u209_u0=~port_687ecc25_;
assign simplePinWrite_u147=and_u935_u0&{1{and_u935_u0}};
assign and_u934_u0=and_u933_u0&and_u945_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3fb682df_u0<=1'h0;
else reg_3fb682df_u0<=and_u935_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_513f5af6_u0<=1'h0;
else reg_513f5af6_u0<=reg_0b0fac36_u0;
end
assign or_u250_u0=reg_513f5af6_result_delayed_u0|and_delayed_u67_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0b0fac36_u0<=1'h0;
else reg_0b0fac36_u0<=reg_3fb682df_result_delayed_u0;
end
assign and_u935_u0=and_u932_u0&and_u945_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u67_u0<=1'h0;
else and_delayed_u67_u0<=and_u934_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3fb682df_result_delayed_u0<=1'h0;
else reg_3fb682df_result_delayed_u0<=reg_3fb682df_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_513f5af6_result_delayed_u0<=1'h0;
else reg_513f5af6_result_delayed_u0<=reg_513f5af6_u0;
end
assign and_u936_u0=and_u944_u0&not_u210_u0;
assign not_u210_u0=~andOp_u96;
assign and_u937_u0=and_u944_u0&andOp_u96;
assign and_u938_u0=and_u943_u0&not_u211_u0;
assign and_u939_u0=and_u943_u0&port_4533a20c_;
assign not_u211_u0=~port_4533a20c_;
assign simplePinWrite_u148=and_u941_u0&{1{and_u941_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4ecbafa0_u0<=1'h0;
else reg_4ecbafa0_u0<=and_delayed_u68_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_78c90025_u0<=1'h0;
else reg_78c90025_u0<=reg_46014afb_u0;
end
assign and_u940_u0=and_u938_u0&and_u943_u0;
assign and_u941_u0=and_u939_u0&and_u943_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u68_u0<=1'h0;
else and_delayed_u68_u0<=and_u941_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_46014afb_u0<=1'h0;
else reg_46014afb_u0<=reg_4ecbafa0_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4ecbafa0_result_delayed_u0<=1'h0;
else reg_4ecbafa0_result_delayed_u0<=reg_4ecbafa0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u69_u0<=1'h0;
else and_delayed_u69_u0<=and_u940_u0;
end
assign or_u251_u0=and_delayed_u69_u0|reg_78c90025_u0;
assign and_u942_u0=and_u936_u0&and_u944_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u70_u0<=1'h0;
else and_delayed_u70_u0<=and_u942_u0;
end
assign or_u252_u0=or_u251_u0|and_delayed_u70_u0;
assign and_u943_u0=and_u937_u0&and_u944_u0;
assign and_u944_u0=and_u931_u0&and_u946_u0;
assign or_u253_u0=and_u935_u0|and_u941_u0;
assign or_u254_u0=or_u250_u0|or_u252_u0;
assign and_u945_u0=and_u930_u0&and_u946_u0;
assign mux_u54_u0=(and_u928_u0)?3'h6:3'h0;
assign or_u255_u0=and_u928_u0|or_u253_u0;
assign and_u946_u0=and_u924_u0&and_u948_u0;
assign or_u256_u0=or_u254_u0|or_u249_u0;
assign and_u947_u0=and_u925_u0&and_u948_u0;
assign or_u257_u0=or_u248_u0|or_u256_u0;
assign and_u948_u0=and_u918_u0&and_u950_u0;
assign mux_u55_u0=(and_u923_u0)?3'h6:{mux_u54_u0[1], mux_u54_u0[1], 1'b0};
assign or_u258_u0=and_u923_u0|or_u255_u0;
assign and_u949_u0=and_u919_u0&and_u950_u0;
assign and_u950_u0=and_u916_u0&and_u717_u0;
assign or_u259_u0=reg_42f13385_u0|or_u257_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_42f13385_u0<=1'h0;
else reg_42f13385_u0<=and_u951_u0;
end
assign and_u951_u0=and_u917_u0&and_u717_u0;
assign midLeftNoConsume2_go_merge=simplePinWrite_u130|simplePinWrite_u142;
assign midLeft2_go_merge=simplePinWrite_u128|simplePinWrite_u140;
assign scoreboard_090d27ac_and=scoreboard_090d27ac_resOr0&scoreboard_090d27ac_resOr1&scoreboard_090d27ac_resOr2&scoreboard_090d27ac_resOr3&scoreboard_090d27ac_resOr4&scoreboard_090d27ac_resOr5;
always @(posedge CLK)
begin
if (bus_07c053e2_)
scoreboard_090d27ac_reg4<=1'h0;
else if (or_u187_u0)
scoreboard_090d27ac_reg4<=1'h1;
else scoreboard_090d27ac_reg4<=scoreboard_090d27ac_reg4;
end
always @(posedge CLK)
begin
if (bus_07c053e2_)
scoreboard_090d27ac_reg0<=1'h0;
else if (or_u229_u0)
scoreboard_090d27ac_reg0<=1'h1;
else scoreboard_090d27ac_reg0<=scoreboard_090d27ac_reg0;
end
always @(posedge CLK)
begin
if (bus_07c053e2_)
scoreboard_090d27ac_reg3<=1'h0;
else if (or_u193_u0)
scoreboard_090d27ac_reg3<=1'h1;
else scoreboard_090d27ac_reg3<=scoreboard_090d27ac_reg3;
end
assign scoreboard_090d27ac_resOr2=or_u205_u0|scoreboard_090d27ac_reg2;
assign scoreboard_090d27ac_resOr0=or_u229_u0|scoreboard_090d27ac_reg0;
always @(posedge CLK)
begin
if (bus_07c053e2_)
scoreboard_090d27ac_reg5<=1'h0;
else if (or_u259_u0)
scoreboard_090d27ac_reg5<=1'h1;
else scoreboard_090d27ac_reg5<=scoreboard_090d27ac_reg5;
end
assign scoreboard_090d27ac_resOr3=or_u193_u0|scoreboard_090d27ac_reg3;
always @(posedge CLK)
begin
if (bus_07c053e2_)
scoreboard_090d27ac_reg2<=1'h0;
else if (or_u205_u0)
scoreboard_090d27ac_reg2<=1'h1;
else scoreboard_090d27ac_reg2<=scoreboard_090d27ac_reg2;
end
assign scoreboard_090d27ac_resOr4=or_u187_u0|scoreboard_090d27ac_reg4;
assign scoreboard_090d27ac_resOr5=or_u259_u0|scoreboard_090d27ac_reg5;
always @(posedge CLK)
begin
if (bus_07c053e2_)
scoreboard_090d27ac_reg1<=1'h0;
else if (or_u247_u0)
scoreboard_090d27ac_reg1<=1'h1;
else scoreboard_090d27ac_reg1<=scoreboard_090d27ac_reg1;
end
assign scoreboard_090d27ac_resOr1=or_u247_u0|scoreboard_090d27ac_reg1;
assign bus_07c053e2_=scoreboard_090d27ac_and|RESET;
assign midLeft1_go_merge=simplePinWrite_u127|simplePinWrite_u139;
assign midLeftNoConsume1_go_merge=simplePinWrite_u129|simplePinWrite_u141;
assign mux_u56_u0=({3{or_u184_u0}}&{2'b0, mux_u44[0]})|({3{and_u734_u0}}&3'h2)|({3{or_u191_u0}}&{2'b1, mux_u45_u0[0]})|({3{or_u204_u0}}&3'h4)|({3{or_u227_u0}}&{2'b10, mux_u49_u0[0]})|({3{or_u246_u0}}&{1'b1, mux_u53_u0[1], 1'b0})|({3{or_u258_u0}}&{mux_u55_u0[1], mux_u55_u0[1], 1'b0});
assign or_u260_u0=or_u184_u0|and_u734_u0|or_u191_u0|or_u204_u0|or_u227_u0|or_u246_u0|or_u258_u0;
assign or_u261_u0=scoreboard_090d27ac_and|reg_12346cc9_result_delayed_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_12346cc9_u0<=1'h0;
else reg_12346cc9_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_12346cc9_result_delayed_u0<=1'h0;
else reg_12346cc9_result_delayed_u0<=reg_12346cc9_u0;
end
assign mux_u57_u0=(GO)?3'h0:mux_u56_u0;
assign or_u262_u0=GO|or_u260_u0;
assign RESULT=or_u262_u0;
assign RESULT_u405=mux_u57_u0;
assign RESULT_u406=simplePinWrite;
assign RESULT_u407=simplePinWrite_u133;
assign RESULT_u408=simplePinWrite_u138;
assign RESULT_u409=simplePinWrite_u144;
assign RESULT_u410=midLeft2_go_merge;
assign RESULT_u411=simplePinWrite_u135;
assign RESULT_u412=simplePinWrite_u143;
assign RESULT_u413=simplePinWrite_u148;
assign RESULT_u414=simplePinWrite_u123;
assign RESULT_u415=simplePinWrite_u137;
assign RESULT_u416=simplePinWrite_u125;
assign RESULT_u417=midLeftNoConsume2_go_merge;
assign RESULT_u418=simplePinWrite_u131;
assign RESULT_u419=simplePinWrite_u147;
assign RESULT_u420=midLeft1_go_merge;
assign RESULT_u421=midLeftNoConsume1_go_merge;
assign RESULT_u422=simplePinWrite_u134;
assign RESULT_u423=simplePinWrite_u126;
assign RESULT_u424=simplePinWrite_u124;
assign RESULT_u425=simplePinWrite_u145;
assign RESULT_u426=simplePinWrite_u136;
assign RESULT_u427=simplePinWrite_u132;
assign RESULT_u428=simplePinWrite_u146;
assign DONE=1'h0;
endmodule



module LL1_L_iunzipFilter2D_bottomLeftNoConsume1(CLK, RESET, GO, port_61b6f9d5_, port_45192321_, port_068d9e17_, port_286032ff_, RESULT, RESULT_u429, RESULT_u430, RESULT_u431, RESULT_u432, RESULT_u433, RESULT_u434, RESULT_u435, RESULT_u436, RESULT_u437, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_61b6f9d5_;
input	[15:0]	port_45192321_;
input		port_068d9e17_;
input	[15:0]	port_286032ff_;
output		RESULT;
output	[15:0]	RESULT_u429;
output		RESULT_u430;
output	[15:0]	RESULT_u431;
output		RESULT_u432;
output	[31:0]	RESULT_u433;
output	[2:0]	RESULT_u434;
output	[15:0]	RESULT_u435;
output	[15:0]	RESULT_u436;
output		RESULT_u437;
output		DONE;
reg		done_cache_u42=1'h0;
wire		and_u952_u0;
wire		or_u263_u0;
reg		done_cache_u43_u0=1'h0;
wire		or_u264_u0;
wire		and_u957_u0;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_3a7bd093_instance_RESULT;
wire	[15:0]	add;
wire	[15:0]	simplePinWrite;
wire		simplePinWrite_u149;
wire	[15:0]	simplePinWrite_u150;
reg		reg_1b5fbf5b_u0=1'h0;
wire		or_u265_u0;
reg		reg_6b4c7d67_u0=1'h0;
reg		reg_51778212_u0=1'h0;
reg		reg_1b5fbf5b_result_delayed_u0=1'h0;
reg		reg_51778212_result_delayed_u0=1'h0;
reg	[15:0]	syncEnable_u31=16'h0;
always @(posedge CLK or posedge GO or posedge or_u263_u0)
begin
if (or_u263_u0)
done_cache_u42<=1'h0;
else if (GO)
done_cache_u42<=1'h1;
else done_cache_u42<=done_cache_u42;
end
assign and_u952_u0=done_cache_u42&port_068d9e17_;
assign or_u263_u0=and_u952_u0|RESET;
always @(posedge CLK or posedge reg_1b5fbf5b_result_delayed_u0 or posedge or_u264_u0)
begin
if (or_u264_u0)
done_cache_u43_u0<=1'h0;
else if (reg_1b5fbf5b_result_delayed_u0)
done_cache_u43_u0<=1'h1;
else done_cache_u43_u0<=done_cache_u43_u0;
end
assign or_u264_u0=and_u957_u0|RESET;
assign and_u957_u0=done_cache_u43_u0&port_068d9e17_;
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_3a7bd093_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_3a7bd093_instance(.GO(reg_51778212_u0), 
  .port_705b5761_(syncEnable_u31), .port_2d505d5c_(port_286032ff_), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_3a7bd093_instance_RESULT));
assign add=port_45192321_+16'h1;
assign simplePinWrite=16'h1&{16{1'h1}};
assign simplePinWrite_u149=reg_51778212_u0&{1{reg_51778212_u0}};
assign simplePinWrite_u150=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_3a7bd093_instance_RESULT&{16{reg_51778212_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1b5fbf5b_u0<=1'h0;
else reg_1b5fbf5b_u0<=GO;
end
assign or_u265_u0=GO|reg_1b5fbf5b_result_delayed_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6b4c7d67_u0<=1'h0;
else reg_6b4c7d67_u0<=reg_51778212_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_51778212_u0<=1'h0;
else reg_51778212_u0<=reg_1b5fbf5b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1b5fbf5b_result_delayed_u0<=1'h0;
else reg_1b5fbf5b_result_delayed_u0<=reg_1b5fbf5b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_51778212_result_delayed_u0<=1'h0;
else reg_51778212_result_delayed_u0<=reg_51778212_u0;
end
always @(posedge CLK)
begin
if (reg_1b5fbf5b_u0)
syncEnable_u31<=port_286032ff_;
end
assign RESULT=GO;
assign RESULT_u429=16'h0;
assign RESULT_u430=GO;
assign RESULT_u431=add;
assign RESULT_u432=or_u265_u0;
assign RESULT_u433=32'h0;
assign RESULT_u434=3'h1;
assign RESULT_u435=simplePinWrite_u150;
assign RESULT_u436=simplePinWrite;
assign RESULT_u437=simplePinWrite_u149;
assign DONE=reg_6b4c7d67_u0;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_3a7bd093_(GO, port_705b5761_, port_2d505d5c_, RESULT);
input		GO;
input	[15:0]	port_705b5761_;
input	[15:0]	port_2d505d5c_;
output	[15:0]	RESULT;
wire	[16:0]	add;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_57123405_instance_RESULT;
assign add={port_705b5761_[15], port_705b5761_}+{port_2d505d5c_[15], port_2d505d5c_};
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_57123405_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_57123405_instance(.GO(GO), 
  .port_01f9e5ba_({add[16], add[16:2]}), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_57123405_instance_RESULT));
assign RESULT=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_57123405_instance_RESULT;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_57123405_(GO, port_01f9e5ba_, RESULT);
input		GO;
input	[15:0]	port_01f9e5ba_;
output	[15:0]	RESULT;
wire		greaterThan;
wire signed	[15:0]	greaterThan_a_signed;
wire signed	[15:0]	greaterThan_b_signed;
wire		and_u961_u0;
wire		and_u962_u0;
wire		not_u212_u0;
wire	[15:0]	mux_u58;
wire		and_u963_u0;
wire		and_u964_u0;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_01f9e5ba_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign and_u961_u0=GO&not_u212_u0;
assign and_u962_u0=GO&greaterThan;
assign not_u212_u0=~greaterThan;
assign mux_u58=(and_u963_u0)?16'h0:port_01f9e5ba_;
assign and_u963_u0=and_u962_u0&GO;
assign and_u964_u0=and_u961_u0&GO;
assign RESULT=mux_u58;
endmodule



module LL1_L_iunzipFilter2D_simplememoryreferee_30774571_(bus_0243864e_, bus_5d3ae11e_, bus_19484e64_, bus_54e8abfe_, bus_20fb712d_, bus_4f73f169_, bus_4279a696_, bus_722d6b97_, bus_1c777956_, bus_13f1caa2_, bus_3bbec1a4_, bus_778a83e5_, bus_21b0d60f_, bus_063abbd4_, bus_2b762ca1_, bus_5dfd93fb_, bus_00516411_, bus_5370ed53_, bus_79564239_, bus_0e3a8226_, bus_04a67cd7_, bus_460823b9_, bus_10bdbe2d_, bus_4a03791e_, bus_51c5155e_, bus_23637f81_, bus_23e6302d_, bus_6eb29e4f_, bus_613d1e04_, bus_5dcadfde_, bus_5c51a8d6_, bus_6767df53_, bus_6fa6325e_, bus_7167efe2_, bus_5884faca_, bus_7b82651c_, bus_12700c62_, bus_78f2c71d_, bus_01cfc67d_, bus_69d0e5eb_, bus_3ae0aed4_, bus_3f2f9d38_, bus_65a9722f_, bus_16b5d3be_, bus_45dfafc9_, bus_35488083_, bus_7f794c6e_, bus_32e4169c_, bus_7247ce17_, bus_3998d8b1_, bus_3df97d91_, bus_5c6c776e_, bus_5ab9a6be_, bus_2d128350_, bus_54e5d40a_, bus_3246468e_, bus_4a5121f7_, bus_5c683fe8_, bus_3189a35f_, bus_1c1d4898_, bus_224fa6f5_, bus_6a39073c_, bus_06490750_, bus_22f52c59_, bus_5ee61a28_, bus_17b97c76_, bus_2346e771_, bus_21b39f31_, bus_15a2faf2_, bus_6ab9c209_, bus_59a547a4_, bus_2eda6c29_, bus_3121b847_, bus_75ed37c9_, bus_7bb56cf6_, bus_577fde87_, bus_0b12336f_, bus_711297cf_, bus_4a8a2bdd_, bus_5968c0b8_, bus_15eaab9b_, bus_14b7951c_, bus_4ab46008_, bus_2f560388_, bus_2e43f4db_, bus_47d6ef03_, bus_1e0f9134_, bus_7f773641_, bus_349b9fac_, bus_3607d9ee_, bus_28bb0475_, bus_170909c9_, bus_4c69ce54_, bus_1ea2aac1_, bus_20897fac_, bus_05cc4bc4_, bus_694f6a4e_, bus_3cc9da1f_, bus_232e245b_, bus_1cb6406c_, bus_7351412b_, bus_45e58a9c_, bus_06fef45c_, bus_1faaec31_, bus_3381d539_, bus_0ca0f630_, bus_317adece_, bus_12ab3e35_, bus_7e595a89_, bus_18c7f89c_, bus_55e3cbdb_, bus_54485535_, bus_4a9b702b_, bus_013fe4a5_, bus_3435fed4_, bus_1ee56c59_, bus_5f8b3986_, bus_59c5b7d5_, bus_2ae9753e_, bus_5a2ebcef_, bus_0ed5862c_, bus_6fff4e52_, bus_4cbd1f1c_, bus_600325c7_, bus_0cb909ae_, bus_62557f73_, bus_42f56b99_, bus_2bae7787_, bus_01a2865d_, bus_5858632d_, bus_516e2378_, bus_34a996e5_);
input		bus_0243864e_;
input		bus_5d3ae11e_;
input		bus_19484e64_;
input	[15:0]	bus_54e8abfe_;
input		bus_20fb712d_;
input		bus_4f73f169_;
input	[15:0]	bus_4279a696_;
input	[31:0]	bus_722d6b97_;
input	[2:0]	bus_1c777956_;
input		bus_13f1caa2_;
input		bus_3bbec1a4_;
input	[15:0]	bus_778a83e5_;
input	[31:0]	bus_21b0d60f_;
input	[2:0]	bus_063abbd4_;
input		bus_2b762ca1_;
input		bus_5dfd93fb_;
input	[15:0]	bus_00516411_;
input	[31:0]	bus_5370ed53_;
input	[2:0]	bus_79564239_;
input		bus_0e3a8226_;
input		bus_04a67cd7_;
input	[15:0]	bus_460823b9_;
input	[31:0]	bus_10bdbe2d_;
input	[2:0]	bus_4a03791e_;
input		bus_51c5155e_;
input		bus_23637f81_;
input	[15:0]	bus_23e6302d_;
input	[31:0]	bus_6eb29e4f_;
input	[2:0]	bus_613d1e04_;
input		bus_5dcadfde_;
input	[31:0]	bus_5c51a8d6_;
input	[2:0]	bus_6767df53_;
input		bus_6fa6325e_;
input	[31:0]	bus_7167efe2_;
input	[2:0]	bus_5884faca_;
input		bus_7b82651c_;
input		bus_12700c62_;
input	[15:0]	bus_78f2c71d_;
input	[31:0]	bus_01cfc67d_;
input	[2:0]	bus_69d0e5eb_;
input		bus_3ae0aed4_;
input		bus_3f2f9d38_;
input	[15:0]	bus_65a9722f_;
input	[31:0]	bus_16b5d3be_;
input	[2:0]	bus_45dfafc9_;
input		bus_35488083_;
input	[31:0]	bus_7f794c6e_;
input	[2:0]	bus_32e4169c_;
input		bus_7247ce17_;
input	[31:0]	bus_3998d8b1_;
input	[2:0]	bus_3df97d91_;
input		bus_5c6c776e_;
input		bus_5ab9a6be_;
input	[15:0]	bus_2d128350_;
input	[31:0]	bus_54e5d40a_;
input	[2:0]	bus_3246468e_;
input		bus_4a5121f7_;
input		bus_5c683fe8_;
input	[15:0]	bus_3189a35f_;
input	[31:0]	bus_1c1d4898_;
input	[2:0]	bus_224fa6f5_;
input		bus_6a39073c_;
input	[31:0]	bus_06490750_;
input	[2:0]	bus_22f52c59_;
input		bus_5ee61a28_;
input	[31:0]	bus_17b97c76_;
input	[2:0]	bus_2346e771_;
input		bus_21b39f31_;
input	[31:0]	bus_15a2faf2_;
input	[2:0]	bus_6ab9c209_;
input		bus_59a547a4_;
input	[31:0]	bus_2eda6c29_;
input	[2:0]	bus_3121b847_;
input		bus_75ed37c9_;
input	[31:0]	bus_7bb56cf6_;
input	[2:0]	bus_577fde87_;
input		bus_0b12336f_;
input	[31:0]	bus_711297cf_;
input	[2:0]	bus_4a8a2bdd_;
input		bus_5968c0b8_;
input	[31:0]	bus_15eaab9b_;
input	[2:0]	bus_14b7951c_;
input		bus_4ab46008_;
input	[31:0]	bus_2f560388_;
input	[2:0]	bus_2e43f4db_;
output	[15:0]	bus_47d6ef03_;
output	[31:0]	bus_1e0f9134_;
output		bus_7f773641_;
output		bus_349b9fac_;
output	[2:0]	bus_3607d9ee_;
output	[15:0]	bus_28bb0475_;
output		bus_170909c9_;
output	[15:0]	bus_4c69ce54_;
output		bus_1ea2aac1_;
output	[15:0]	bus_20897fac_;
output		bus_05cc4bc4_;
output	[15:0]	bus_694f6a4e_;
output		bus_3cc9da1f_;
output	[15:0]	bus_232e245b_;
output		bus_1cb6406c_;
output	[15:0]	bus_7351412b_;
output		bus_45e58a9c_;
output	[15:0]	bus_06fef45c_;
output		bus_1faaec31_;
output	[15:0]	bus_3381d539_;
output		bus_0ca0f630_;
output	[15:0]	bus_317adece_;
output		bus_12ab3e35_;
output	[15:0]	bus_7e595a89_;
output		bus_18c7f89c_;
output	[15:0]	bus_55e3cbdb_;
output		bus_54485535_;
output	[15:0]	bus_4a9b702b_;
output		bus_013fe4a5_;
output	[15:0]	bus_3435fed4_;
output		bus_1ee56c59_;
output	[15:0]	bus_5f8b3986_;
output		bus_59c5b7d5_;
output	[15:0]	bus_2ae9753e_;
output		bus_5a2ebcef_;
output	[15:0]	bus_0ed5862c_;
output		bus_6fff4e52_;
output	[15:0]	bus_4cbd1f1c_;
output		bus_600325c7_;
output	[15:0]	bus_0cb909ae_;
output		bus_62557f73_;
output	[15:0]	bus_42f56b99_;
output		bus_2bae7787_;
output	[15:0]	bus_01a2865d_;
output		bus_5858632d_;
output	[15:0]	bus_516e2378_;
output		bus_34a996e5_;
reg		done_qual_u21=1'h0;
wire		and_48004704_u0;
wire		not_0f03d606_u0;
reg		done_qual_u22_u0=1'h0;
reg		done_qual_u23_u0=1'h0;
wire		not_57294c3d_u0;
reg		done_qual_u24_u0=1'h0;
wire		or_61c9d2d2_u0;
wire		and_744ff554_u0;
wire		and_1d963f8b_u0;
wire	[15:0]	mux_386b5075_u0;
wire		or_443ea220_u0;
wire		not_0fd3facd_u0;
wire		not_0e02b922_u0;
wire		or_376ca44e_u0;
reg		done_qual_u25_u0=1'h0;
reg		done_qual_u26_u0=1'h0;
reg		done_qual_u27_u0=1'h0;
reg		done_qual_u28_u0=1'h0;
wire		not_5d9b3eb0_u0;
wire		or_42446b6a_u0;
wire		not_3fb04681_u0;
wire		or_68322601_u0;
wire		or_4f58176b_u0;
wire		or_6e7b574e_u0;
reg		done_qual_u29_u0=1'h0;
wire		not_6121231a_u0;
wire		and_558cbac8_u0;
reg		done_qual_u30_u0=1'h0;
wire		and_35034448_u0;
wire		not_652f977e_u0;
wire		or_49525606_u0;
wire		or_47221076_u0;
wire		or_632b937d_u0;
wire		or_05b67fed_u0;
wire		not_4e329d6c_u0;
reg		done_qual_u31_u0=1'h0;
reg		done_qual_u32_u0=1'h0;
wire		and_2ca435c1_u0;
wire		not_0ae43781_u0;
wire		and_0596a1fe_u0;
wire		or_15a77fcd_u0;
reg		done_qual_u33_u0=1'h0;
reg		done_qual_u34_u0=1'h0;
wire		or_5a58e728_u0;
wire		or_08831bf3_u0;
wire		and_03c397b1_u0;
wire		not_129bafe9_u0;
wire		not_208a2ef0_u0;
wire		and_36952de9_u0;
wire		and_46cceeb2_u0;
wire		not_265b09db_u0;
reg		done_qual_u35_u0=1'h0;
wire		or_73d64a57_u0;
wire		and_366a77e8_u0;
wire		and_434102c7_u0;
wire		or_28a78e20_u0;
wire		or_6fe1506a_u0;
wire		and_34a50537_u0;
wire		or_141acb8e_u0;
wire		or_34f53461_u0;
wire		or_0990f908_u0;
wire		and_222709be_u0;
wire		not_66b88021_u0;
wire		or_48fb5867_u0;
reg		done_qual_u36_u0=1'h0;
wire		not_075daac2_u0;
wire	[31:0]	mux_5955d3f5_u0;
wire		not_7b6d03cd_u0;
wire		or_4c5da1fc_u0;
wire		or_02c9dc66_u0;
wire		not_63307580_u0;
reg		done_qual_u37_u0=1'h0;
reg		done_qual_u38_u0=1'h0;
wire		or_0ac6677a_u0;
wire		or_5cdcdf63_u0;
wire		or_1a61a0a0_u0;
wire		and_1fac886f_u0;
wire		and_44bc7676_u0;
wire		not_11fe5934_u0;
wire		and_0578f3ae_u0;
wire		or_2767e7bd_u0;
reg		done_qual_u39_u0=1'h0;
wire		and_6e3d1cdf_u0;
reg		done_qual_u40_u0=1'h0;
wire		and_08ad8d45_u0;
wire		not_541640ff_u0;
reg		done_qual_u41_u0=1'h0;
wire		not_50bfcb55_u0;
wire		and_71e11313_u0;
wire		and_2f0bb9f9_u0;
wire		or_3f943b60_u0;
wire		or_4b83ad74_u0;
wire		or_74b2564b_u0;
wire		not_320ffcf5_u0;
wire		or_27bb9f44_u0;
wire		or_310ea7f1_u0;
always @(posedge bus_0243864e_)
begin
if (bus_5d3ae11e_)
done_qual_u21<=1'h0;
else done_qual_u21<=bus_6a39073c_;
end
assign and_48004704_u0=or_15a77fcd_u0&bus_19484e64_;
assign not_0f03d606_u0=~bus_19484e64_;
always @(posedge bus_0243864e_)
begin
if (bus_5d3ae11e_)
done_qual_u22_u0<=1'h0;
else done_qual_u22_u0<=or_5cdcdf63_u0;
end
always @(posedge bus_0243864e_)
begin
if (bus_5d3ae11e_)
done_qual_u23_u0<=1'h0;
else done_qual_u23_u0<=or_08831bf3_u0;
end
assign not_57294c3d_u0=~bus_19484e64_;
always @(posedge bus_0243864e_)
begin
if (bus_5d3ae11e_)
done_qual_u24_u0<=1'h0;
else done_qual_u24_u0<=bus_6fa6325e_;
end
assign or_61c9d2d2_u0=or_49525606_u0|done_qual_u41_u0;
assign and_744ff554_u0=or_2767e7bd_u0&bus_19484e64_;
assign and_1d963f8b_u0=or_4f58176b_u0&bus_19484e64_;
assign mux_386b5075_u0=({16{bus_4f73f169_}}&bus_4279a696_)|({16{bus_3bbec1a4_}}&bus_778a83e5_)|({16{bus_5dfd93fb_}}&bus_00516411_)|({16{bus_04a67cd7_}}&bus_460823b9_)|({16{bus_23637f81_}}&bus_23e6302d_)|({16{bus_12700c62_}}&bus_78f2c71d_)|({16{bus_3f2f9d38_}}&bus_65a9722f_)|({16{bus_5ab9a6be_}}&bus_2d128350_)|({16{bus_5c683fe8_}}&bus_3189a35f_);
assign or_443ea220_u0=bus_2b762ca1_|bus_5dfd93fb_;
assign not_0fd3facd_u0=~bus_19484e64_;
assign not_0e02b922_u0=~bus_19484e64_;
assign or_376ca44e_u0=bus_4a5121f7_|bus_5c683fe8_;
always @(posedge bus_0243864e_)
begin
if (bus_5d3ae11e_)
done_qual_u25_u0<=1'h0;
else done_qual_u25_u0<=bus_21b39f31_;
end
always @(posedge bus_0243864e_)
begin
if (bus_5d3ae11e_)
done_qual_u26_u0<=1'h0;
else done_qual_u26_u0<=bus_5968c0b8_;
end
always @(posedge bus_0243864e_)
begin
if (bus_5d3ae11e_)
done_qual_u27_u0<=1'h0;
else done_qual_u27_u0<=or_310ea7f1_u0;
end
always @(posedge bus_0243864e_)
begin
if (bus_5d3ae11e_)
done_qual_u28_u0<=1'h0;
else done_qual_u28_u0<=bus_5ee61a28_;
end
assign not_5d9b3eb0_u0=~bus_19484e64_;
assign or_42446b6a_u0=bus_59a547a4_|done_qual_u33_u0;
assign not_3fb04681_u0=~bus_19484e64_;
assign or_68322601_u0=or_5cdcdf63_u0|done_qual_u22_u0;
assign or_4f58176b_u0=bus_75ed37c9_|done_qual_u31_u0;
assign or_6e7b574e_u0=bus_5968c0b8_|done_qual_u26_u0;
always @(posedge bus_0243864e_)
begin
if (bus_5d3ae11e_)
done_qual_u29_u0<=1'h0;
else done_qual_u29_u0<=or_443ea220_u0;
end
assign not_6121231a_u0=~bus_19484e64_;
assign and_558cbac8_u0=or_28a78e20_u0&bus_19484e64_;
always @(posedge bus_0243864e_)
begin
if (bus_5d3ae11e_)
done_qual_u30_u0<=1'h0;
else done_qual_u30_u0<=bus_7247ce17_;
end
assign and_35034448_u0=or_0990f908_u0&bus_19484e64_;
assign not_652f977e_u0=~bus_19484e64_;
assign or_49525606_u0=bus_20fb712d_|bus_4f73f169_;
assign or_47221076_u0=or_141acb8e_u0|done_qual_u35_u0;
assign or_632b937d_u0=or_376ca44e_u0|done_qual_u39_u0;
assign or_05b67fed_u0=bus_7b82651c_|bus_12700c62_;
assign not_4e329d6c_u0=~bus_19484e64_;
always @(posedge bus_0243864e_)
begin
if (bus_5d3ae11e_)
done_qual_u31_u0<=1'h0;
else done_qual_u31_u0<=bus_75ed37c9_;
end
always @(posedge bus_0243864e_)
begin
if (bus_5d3ae11e_)
done_qual_u32_u0<=1'h0;
else done_qual_u32_u0<=bus_0b12336f_;
end
assign and_2ca435c1_u0=or_27bb9f44_u0&bus_19484e64_;
assign not_0ae43781_u0=~bus_19484e64_;
assign and_0596a1fe_u0=or_632b937d_u0&bus_19484e64_;
assign or_15a77fcd_u0=or_443ea220_u0|done_qual_u29_u0;
always @(posedge bus_0243864e_)
begin
if (bus_5d3ae11e_)
done_qual_u33_u0<=1'h0;
else done_qual_u33_u0<=bus_59a547a4_;
end
always @(posedge bus_0243864e_)
begin
if (bus_5d3ae11e_)
done_qual_u34_u0<=1'h0;
else done_qual_u34_u0<=bus_4ab46008_;
end
assign or_5a58e728_u0=or_49525606_u0|or_5cdcdf63_u0|or_443ea220_u0|or_08831bf3_u0|or_141acb8e_u0|bus_5dcadfde_|bus_6fa6325e_|or_05b67fed_u0|or_34f53461_u0|bus_35488083_|bus_7247ce17_|or_310ea7f1_u0|or_376ca44e_u0|bus_6a39073c_|bus_5ee61a28_|bus_21b39f31_|bus_59a547a4_|bus_75ed37c9_|bus_0b12336f_|bus_5968c0b8_|bus_4ab46008_;
assign or_08831bf3_u0=bus_0e3a8226_|bus_04a67cd7_;
assign and_03c397b1_u0=or_68322601_u0&bus_19484e64_;
assign not_129bafe9_u0=~bus_19484e64_;
assign not_208a2ef0_u0=~bus_19484e64_;
assign and_36952de9_u0=or_47221076_u0&bus_19484e64_;
assign and_46cceeb2_u0=or_48fb5867_u0&bus_19484e64_;
assign not_265b09db_u0=~bus_19484e64_;
always @(posedge bus_0243864e_)
begin
if (bus_5d3ae11e_)
done_qual_u35_u0<=1'h0;
else done_qual_u35_u0<=or_141acb8e_u0;
end
assign or_73d64a57_u0=bus_0b12336f_|done_qual_u32_u0;
assign and_366a77e8_u0=or_1a61a0a0_u0&bus_19484e64_;
assign and_434102c7_u0=or_42446b6a_u0&bus_19484e64_;
assign or_28a78e20_u0=bus_7247ce17_|done_qual_u30_u0;
assign or_6fe1506a_u0=or_08831bf3_u0|done_qual_u23_u0;
assign and_34a50537_u0=or_02c9dc66_u0&bus_19484e64_;
assign or_141acb8e_u0=bus_51c5155e_|bus_23637f81_;
assign or_34f53461_u0=bus_3ae0aed4_|bus_3f2f9d38_;
assign or_0990f908_u0=bus_21b39f31_|done_qual_u25_u0;
assign and_222709be_u0=or_61c9d2d2_u0&bus_19484e64_;
assign not_66b88021_u0=~bus_19484e64_;
assign or_48fb5867_u0=bus_4ab46008_|done_qual_u34_u0;
assign bus_47d6ef03_=mux_386b5075_u0;
assign bus_1e0f9134_=mux_5955d3f5_u0;
assign bus_7f773641_=or_3f943b60_u0;
assign bus_349b9fac_=or_5a58e728_u0;
assign bus_3607d9ee_=3'h1;
assign bus_28bb0475_=bus_54e8abfe_;
assign bus_170909c9_=and_222709be_u0;
assign bus_4c69ce54_=bus_54e8abfe_;
assign bus_1ea2aac1_=and_03c397b1_u0;
assign bus_20897fac_=bus_54e8abfe_;
assign bus_05cc4bc4_=and_48004704_u0;
assign bus_694f6a4e_=bus_54e8abfe_;
assign bus_3cc9da1f_=and_71e11313_u0;
assign bus_232e245b_=bus_54e8abfe_;
assign bus_1cb6406c_=and_36952de9_u0;
assign bus_7351412b_=bus_54e8abfe_;
assign bus_45e58a9c_=and_366a77e8_u0;
assign bus_06fef45c_=bus_54e8abfe_;
assign bus_1faaec31_=and_44bc7676_u0;
assign bus_3381d539_=bus_54e8abfe_;
assign bus_0ca0f630_=and_34a50537_u0;
assign bus_317adece_=bus_54e8abfe_;
assign bus_12ab3e35_=and_2f0bb9f9_u0;
assign bus_7e595a89_=bus_54e8abfe_;
assign bus_18c7f89c_=and_2ca435c1_u0;
assign bus_55e3cbdb_=bus_54e8abfe_;
assign bus_54485535_=and_558cbac8_u0;
assign bus_4a9b702b_=bus_54e8abfe_;
assign bus_013fe4a5_=and_1fac886f_u0;
assign bus_3435fed4_=bus_54e8abfe_;
assign bus_1ee56c59_=and_0596a1fe_u0;
assign bus_5f8b3986_=bus_54e8abfe_;
assign bus_59c5b7d5_=and_744ff554_u0;
assign bus_2ae9753e_=bus_54e8abfe_;
assign bus_5a2ebcef_=and_0578f3ae_u0;
assign bus_0ed5862c_=bus_54e8abfe_;
assign bus_6fff4e52_=and_35034448_u0;
assign bus_4cbd1f1c_=bus_54e8abfe_;
assign bus_600325c7_=and_434102c7_u0;
assign bus_0cb909ae_=bus_54e8abfe_;
assign bus_62557f73_=and_1d963f8b_u0;
assign bus_42f56b99_=bus_54e8abfe_;
assign bus_2bae7787_=and_6e3d1cdf_u0;
assign bus_01a2865d_=bus_54e8abfe_;
assign bus_5858632d_=and_08ad8d45_u0;
assign bus_516e2378_=bus_54e8abfe_;
assign bus_34a996e5_=and_46cceeb2_u0;
always @(posedge bus_0243864e_)
begin
if (bus_5d3ae11e_)
done_qual_u36_u0<=1'h0;
else done_qual_u36_u0<=bus_5dcadfde_;
end
assign not_075daac2_u0=~bus_19484e64_;
assign mux_5955d3f5_u0=({32{or_49525606_u0}}&bus_722d6b97_)|({32{or_5cdcdf63_u0}}&32'h0)|({32{or_443ea220_u0}}&32'h0)|({32{or_08831bf3_u0}}&32'h0)|({32{or_141acb8e_u0}}&32'h0)|({32{bus_5dcadfde_}}&32'h0)|({32{bus_6fa6325e_}}&32'h0)|({32{or_05b67fed_u0}}&32'h0)|({32{or_34f53461_u0}}&32'h0)|({32{bus_35488083_}}&32'h0)|({32{bus_7247ce17_}}&32'h0)|({32{or_310ea7f1_u0}}&32'h0)|({32{or_376ca44e_u0}}&32'h0)|({32{bus_6a39073c_}}&32'h0)|({32{bus_5ee61a28_}}&32'h0)|({32{bus_21b39f31_}}&32'h0)|({32{bus_59a547a4_}}&32'h0)|({32{bus_75ed37c9_}}&32'h0)|({32{bus_0b12336f_}}&32'h0)|({32{bus_5968c0b8_}}&32'h0)|({32{bus_4ab46008_}}&32'h0);
assign not_7b6d03cd_u0=~bus_19484e64_;
assign or_4c5da1fc_u0=bus_6fa6325e_|done_qual_u24_u0;
assign or_02c9dc66_u0=or_05b67fed_u0|done_qual_u40_u0;
assign not_63307580_u0=~bus_19484e64_;
always @(posedge bus_0243864e_)
begin
if (bus_5d3ae11e_)
done_qual_u37_u0<=1'h0;
else done_qual_u37_u0<=bus_35488083_;
end
always @(posedge bus_0243864e_)
begin
if (bus_5d3ae11e_)
done_qual_u38_u0<=1'h0;
else done_qual_u38_u0<=or_34f53461_u0;
end
assign or_0ac6677a_u0=bus_5ee61a28_|done_qual_u28_u0;
assign or_5cdcdf63_u0=bus_13f1caa2_|bus_3bbec1a4_;
assign or_1a61a0a0_u0=bus_5dcadfde_|done_qual_u36_u0;
assign and_1fac886f_u0=or_4b83ad74_u0&bus_19484e64_;
assign and_44bc7676_u0=or_4c5da1fc_u0&bus_19484e64_;
assign not_11fe5934_u0=~bus_19484e64_;
assign and_0578f3ae_u0=or_0ac6677a_u0&bus_19484e64_;
assign or_2767e7bd_u0=bus_6a39073c_|done_qual_u21;
always @(posedge bus_0243864e_)
begin
if (bus_5d3ae11e_)
done_qual_u39_u0<=1'h0;
else done_qual_u39_u0<=or_376ca44e_u0;
end
assign and_6e3d1cdf_u0=or_73d64a57_u0&bus_19484e64_;
always @(posedge bus_0243864e_)
begin
if (bus_5d3ae11e_)
done_qual_u40_u0<=1'h0;
else done_qual_u40_u0<=or_05b67fed_u0;
end
assign and_08ad8d45_u0=or_6e7b574e_u0&bus_19484e64_;
assign not_541640ff_u0=~bus_19484e64_;
always @(posedge bus_0243864e_)
begin
if (bus_5d3ae11e_)
done_qual_u41_u0<=1'h0;
else done_qual_u41_u0<=or_49525606_u0;
end
assign not_50bfcb55_u0=~bus_19484e64_;
assign and_71e11313_u0=or_6fe1506a_u0&bus_19484e64_;
assign and_2f0bb9f9_u0=or_74b2564b_u0&bus_19484e64_;
assign or_3f943b60_u0=bus_4f73f169_|bus_3bbec1a4_|bus_5dfd93fb_|bus_04a67cd7_|bus_23637f81_|bus_12700c62_|bus_3f2f9d38_|bus_5ab9a6be_|bus_5c683fe8_;
assign or_4b83ad74_u0=or_310ea7f1_u0|done_qual_u27_u0;
assign or_74b2564b_u0=or_34f53461_u0|done_qual_u38_u0;
assign not_320ffcf5_u0=~bus_19484e64_;
assign or_27bb9f44_u0=bus_35488083_|done_qual_u37_u0;
assign or_310ea7f1_u0=bus_5c6c776e_|bus_5ab9a6be_;
endmodule



module LL1_L_iunzipFilter2D_topRight(CLK, RESET, GO, port_441cd972_, port_7fcde167_, port_05ea2457_, port_6215fb35_, port_4a4dafea_, port_50ff8e8d_, RESULT, RESULT_u438, RESULT_u439, RESULT_u440, RESULT_u441, RESULT_u442, RESULT_u443, RESULT_u444, RESULT_u445, RESULT_u446, RESULT_u447, RESULT_u448, RESULT_u449, RESULT_u450, RESULT_u451, RESULT_u452, RESULT_u453, RESULT_u454, RESULT_u455, RESULT_u456, RESULT_u457, DONE);
input		CLK;
input		RESET;
input		GO;
input	[31:0]	port_441cd972_;
input		port_7fcde167_;
input		port_05ea2457_;
input	[15:0]	port_6215fb35_;
input		port_4a4dafea_;
input	[15:0]	port_50ff8e8d_;
output		RESULT;
output	[31:0]	RESULT_u438;
output		RESULT_u439;
output	[15:0]	RESULT_u440;
output		RESULT_u441;
output	[15:0]	RESULT_u442;
output		RESULT_u443;
output	[15:0]	RESULT_u444;
output		RESULT_u445;
output		RESULT_u446;
output		RESULT_u447;
output	[31:0]	RESULT_u448;
output	[2:0]	RESULT_u449;
output		RESULT_u450;
output	[31:0]	RESULT_u451;
output	[15:0]	RESULT_u452;
output	[2:0]	RESULT_u453;
output	[15:0]	RESULT_u454;
output	[15:0]	RESULT_u455;
output		RESULT_u456;
output		RESULT_u457;
output		DONE;
wire		simplePinWrite;
wire		or_u266_u0;
reg		done_cache_u44=1'h0;
wire		and_u967_u0;
wire		and_u971_u0;
reg		done_cache_u45_u0=1'h0;
wire		or_u267_u0;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_1d713b85_instance_RESULT;
wire		or_u268_u0;
reg		reg_62c182f7_u0=1'h0;
wire		and_u980_u0;
wire	[31:0]	add;
wire		not_u214;
wire	[15:0]	simplePinWrite_u151;
wire	[15:0]	simplePinWrite_u152;
wire		simplePinWrite_u153;
reg		reg_4ad734d1_u0=1'h0;
reg	[15:0]	syncEnable_u32=16'h0;
reg	[15:0]	syncEnable_u33_u0=16'h0;
reg		reg_53c0809f_u0=1'h0;
reg		reg_749d0fe6_u0=1'h0;
reg		reg_749d0fe6_result_delayed_u0=1'h0;
wire		or_u269_u0;
reg		reg_4ad734d1_result_delayed_u0=1'h0;
reg		reg_4ad734d1_result_delayed_result_delayed_u0=1'h0;
assign simplePinWrite=GO&{1{GO}};
assign or_u266_u0=and_u967_u0|RESET;
always @(posedge CLK or posedge GO or posedge or_u266_u0)
begin
if (or_u266_u0)
done_cache_u44<=1'h0;
else if (GO)
done_cache_u44<=1'h1;
else done_cache_u44<=done_cache_u44;
end
assign and_u967_u0=done_cache_u44&port_4a4dafea_;
assign and_u971_u0=done_cache_u45_u0&port_4a4dafea_;
always @(posedge CLK or posedge reg_749d0fe6_result_delayed_u0 or posedge or_u267_u0)
begin
if (or_u267_u0)
done_cache_u45_u0<=1'h0;
else if (reg_749d0fe6_result_delayed_u0)
done_cache_u45_u0<=1'h1;
else done_cache_u45_u0<=done_cache_u45_u0;
end
assign or_u267_u0=and_u971_u0|RESET;
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_1d713b85_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_1d713b85_instance(.GO(reg_53c0809f_u0), 
  .port_69b16870_(port_6215fb35_), .port_0216e718_(syncEnable_u32), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_1d713b85_instance_RESULT));
assign or_u268_u0=and_u980_u0|RESET;
always @(posedge CLK or posedge reg_4ad734d1_result_delayed_u0 or posedge or_u268_u0)
begin
if (or_u268_u0)
reg_62c182f7_u0<=1'h0;
else if (reg_4ad734d1_result_delayed_u0)
reg_62c182f7_u0<=1'h1;
else reg_62c182f7_u0<=reg_62c182f7_u0;
end
assign and_u980_u0=reg_62c182f7_u0&port_4a4dafea_;
assign add=port_441cd972_+32'h1;
assign not_u214=!port_7fcde167_;
assign simplePinWrite_u151=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_1d713b85_instance_RESULT&{16{reg_53c0809f_u0}};
assign simplePinWrite_u152=16'h1&{16{1'h1}};
assign simplePinWrite_u153=reg_53c0809f_u0&{1{reg_53c0809f_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4ad734d1_u0<=1'h0;
else reg_4ad734d1_u0<=reg_53c0809f_u0;
end
always @(posedge CLK)
begin
if (reg_749d0fe6_u0)
syncEnable_u32<=port_6215fb35_;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u33_u0<=port_50ff8e8d_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_53c0809f_u0<=1'h0;
else reg_53c0809f_u0<=reg_749d0fe6_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_749d0fe6_u0<=1'h0;
else reg_749d0fe6_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_749d0fe6_result_delayed_u0<=1'h0;
else reg_749d0fe6_result_delayed_u0<=reg_749d0fe6_u0;
end
assign or_u269_u0=GO|reg_749d0fe6_result_delayed_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4ad734d1_result_delayed_u0<=1'h0;
else reg_4ad734d1_result_delayed_u0<=reg_4ad734d1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4ad734d1_result_delayed_result_delayed_u0<=1'h0;
else reg_4ad734d1_result_delayed_result_delayed_u0<=reg_4ad734d1_result_delayed_u0;
end
assign RESULT=GO;
assign RESULT_u438=add;
assign RESULT_u439=GO;
assign RESULT_u440=16'h0;
assign RESULT_u441=GO;
assign RESULT_u442=16'h0;
assign RESULT_u443=GO;
assign RESULT_u444=16'h1;
assign RESULT_u445=GO;
assign RESULT_u446=not_u214;
assign RESULT_u447=or_u269_u0;
assign RESULT_u448=32'h0;
assign RESULT_u449=3'h1;
assign RESULT_u450=reg_4ad734d1_result_delayed_u0;
assign RESULT_u451=32'h0;
assign RESULT_u452=syncEnable_u33_u0;
assign RESULT_u453=3'h1;
assign RESULT_u454=simplePinWrite_u151;
assign RESULT_u455=simplePinWrite_u152;
assign RESULT_u456=simplePinWrite;
assign RESULT_u457=simplePinWrite_u153;
assign DONE=reg_4ad734d1_result_delayed_result_delayed_u0;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_1d713b85_(GO, port_69b16870_, port_0216e718_, RESULT);
input		GO;
input	[15:0]	port_69b16870_;
input	[15:0]	port_0216e718_;
output	[15:0]	RESULT;
wire	[16:0]	add;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_364c9329_instance_RESULT;
assign add={port_0216e718_[15], port_0216e718_}+{port_69b16870_[15], port_69b16870_};
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_364c9329_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_364c9329_instance(.GO(GO), 
  .port_38957502_({add[16], add[16:2]}), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_364c9329_instance_RESULT));
assign RESULT=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_364c9329_instance_RESULT;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_364c9329_(GO, port_38957502_, RESULT);
input		GO;
input	[15:0]	port_38957502_;
output	[15:0]	RESULT;
wire		greaterThan;
wire signed	[15:0]	greaterThan_a_signed;
wire signed	[15:0]	greaterThan_b_signed;
wire		and_u975_u0;
wire		and_u976_u0;
wire		not_u213_u0;
wire		and_u977_u0;
wire	[15:0]	mux_u59;
wire		and_u978_u0;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_38957502_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign and_u975_u0=GO&not_u213_u0;
assign and_u976_u0=GO&greaterThan;
assign not_u213_u0=~greaterThan;
assign and_u977_u0=and_u976_u0&GO;
assign mux_u59=(and_u977_u0)?16'h0:port_38957502_;
assign and_u978_u0=and_u975_u0&GO;
assign RESULT=mux_u59;
endmodule



module LL1_L_iunzipFilter2D_globalreset_physical_3810141d_(bus_3dc23f78_, bus_2f4fdc33_, bus_7290ab84_);
input		bus_3dc23f78_;
input		bus_2f4fdc33_;
output		bus_7290ab84_;
reg		glitch_u13=1'h0;
wire		or_6e19f5bb_u0;
wire		not_25c2c281_u0;
reg		sample_u13=1'h0;
wire		and_79251d79_u0;
reg		final_u13=1'h1;
reg		cross_u13=1'h0;
always @(posedge bus_3dc23f78_)
begin
glitch_u13<=cross_u13;
end
assign or_6e19f5bb_u0=bus_2f4fdc33_|final_u13;
assign not_25c2c281_u0=~and_79251d79_u0;
assign bus_7290ab84_=or_6e19f5bb_u0;
always @(posedge bus_3dc23f78_)
begin
sample_u13<=1'h1;
end
assign and_79251d79_u0=cross_u13&glitch_u13;
always @(posedge bus_3dc23f78_)
begin
final_u13<=not_25c2c281_u0;
end
always @(posedge bus_3dc23f78_)
begin
cross_u13<=sample_u13;
end
endmodule



module LL1_L_iunzipFilter2D_midLeft2(CLK, RESET, GO, port_38ad9985_, port_56487516_, port_17d61741_, port_0d7c2f45_, port_43399a57_, port_58424af2_, port_541437a9_, RESULT, RESULT_u458, RESULT_u459, RESULT_u460, RESULT_u461, RESULT_u462, RESULT_u463, RESULT_u464, RESULT_u465, RESULT_u466, RESULT_u467, RESULT_u468, RESULT_u469, RESULT_u470, RESULT_u471, RESULT_u472, RESULT_u473, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_38ad9985_;
input	[31:0]	port_56487516_;
input	[15:0]	port_17d61741_;
input		port_0d7c2f45_;
input	[15:0]	port_43399a57_;
input		port_58424af2_;
input	[15:0]	port_541437a9_;
output		RESULT;
output	[15:0]	RESULT_u458;
output		RESULT_u459;
output	[31:0]	RESULT_u460;
output		RESULT_u461;
output	[15:0]	RESULT_u462;
output		RESULT_u463;
output	[31:0]	RESULT_u464;
output	[2:0]	RESULT_u465;
output		RESULT_u466;
output	[31:0]	RESULT_u467;
output	[15:0]	RESULT_u468;
output	[2:0]	RESULT_u469;
output	[15:0]	RESULT_u470;
output		RESULT_u471;
output	[15:0]	RESULT_u472;
output		RESULT_u473;
output		DONE;
wire		simplePinWrite;
wire		and_u982_u0;
wire		or_u270_u0;
reg		done_cache_u46=1'h0;
wire		or_u271_u0;
reg		done_cache_u47_u0=1'h0;
wire		and_u987_u0;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_1568113c_instance_RESULT;
wire		or_u272_u0;
reg		reg_116e9bd8_u0=1'h0;
wire		and_u996_u0;
wire	[31:0]	add;
wire	[15:0]	add_u12;
wire	[15:0]	simplePinWrite_u154;
wire	[15:0]	simplePinWrite_u155;
wire		simplePinWrite_u156;
reg	[15:0]	syncEnable_u34=16'h0;
reg		reg_3dea818b_u0=1'h0;
reg	[15:0]	syncEnable_u35_u0=16'h0;
wire		or_u273_u0;
reg		reg_36b3f317_u0=1'h0;
reg		reg_5d4c5781_u0=1'h0;
reg		reg_2761b2b1_u0=1'h0;
reg		reg_36b3f317_result_delayed_u0=1'h0;
reg		reg_3dea818b_result_delayed_u0=1'h0;
assign simplePinWrite=GO&{1{GO}};
assign and_u982_u0=done_cache_u46&port_58424af2_;
assign or_u270_u0=and_u982_u0|RESET;
always @(posedge CLK or posedge GO or posedge or_u270_u0)
begin
if (or_u270_u0)
done_cache_u46<=1'h0;
else if (GO)
done_cache_u46<=1'h1;
else done_cache_u46<=done_cache_u46;
end
assign or_u271_u0=and_u987_u0|RESET;
always @(posedge CLK or posedge reg_5d4c5781_u0 or posedge or_u271_u0)
begin
if (or_u271_u0)
done_cache_u47_u0<=1'h0;
else if (reg_5d4c5781_u0)
done_cache_u47_u0<=1'h1;
else done_cache_u47_u0<=done_cache_u47_u0;
end
assign and_u987_u0=done_cache_u47_u0&port_58424af2_;
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_1568113c_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_1568113c_instance(.GO(reg_36b3f317_u0), 
  .port_4553943c_(syncEnable_u35_u0), .port_5a6712aa_(port_43399a57_), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_1568113c_instance_RESULT));
assign or_u272_u0=and_u996_u0|RESET;
always @(posedge CLK or posedge reg_3dea818b_u0 or posedge or_u272_u0)
begin
if (or_u272_u0)
reg_116e9bd8_u0<=1'h0;
else if (reg_3dea818b_u0)
reg_116e9bd8_u0<=1'h1;
else reg_116e9bd8_u0<=reg_116e9bd8_u0;
end
assign and_u996_u0=reg_116e9bd8_u0&port_58424af2_;
assign add=port_56487516_+32'h1;
assign add_u12=port_17d61741_+16'h1;
assign simplePinWrite_u154=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_1568113c_instance_RESULT&{16{reg_36b3f317_u0}};
assign simplePinWrite_u155=16'h1&{16{1'h1}};
assign simplePinWrite_u156=reg_36b3f317_u0&{1{reg_36b3f317_u0}};
always @(posedge CLK)
begin
if (GO)
syncEnable_u34<=port_541437a9_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3dea818b_u0<=1'h0;
else reg_3dea818b_u0<=reg_36b3f317_result_delayed_u0;
end
always @(posedge CLK)
begin
if (reg_2761b2b1_u0)
syncEnable_u35_u0<=port_43399a57_;
end
assign or_u273_u0=GO|reg_5d4c5781_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_36b3f317_u0<=1'h0;
else reg_36b3f317_u0<=reg_5d4c5781_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5d4c5781_u0<=1'h0;
else reg_5d4c5781_u0<=reg_2761b2b1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2761b2b1_u0<=1'h0;
else reg_2761b2b1_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_36b3f317_result_delayed_u0<=1'h0;
else reg_36b3f317_result_delayed_u0<=reg_36b3f317_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3dea818b_result_delayed_u0<=1'h0;
else reg_3dea818b_result_delayed_u0<=reg_3dea818b_u0;
end
assign RESULT=GO;
assign RESULT_u458=16'h0;
assign RESULT_u459=GO;
assign RESULT_u460=add;
assign RESULT_u461=GO;
assign RESULT_u462=add_u12;
assign RESULT_u463=or_u273_u0;
assign RESULT_u464=32'h0;
assign RESULT_u465=3'h1;
assign RESULT_u466=reg_3dea818b_u0;
assign RESULT_u467=32'h0;
assign RESULT_u468=syncEnable_u34;
assign RESULT_u469=3'h1;
assign RESULT_u470=simplePinWrite_u154;
assign RESULT_u471=simplePinWrite;
assign RESULT_u472=simplePinWrite_u155;
assign RESULT_u473=simplePinWrite_u156;
assign DONE=reg_3dea818b_result_delayed_u0;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_1568113c_(GO, port_4553943c_, port_5a6712aa_, RESULT);
input		GO;
input	[15:0]	port_4553943c_;
input	[15:0]	port_5a6712aa_;
output	[15:0]	RESULT;
wire	[15:0]	subtract;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_5d300b1c_instance_RESULT;
assign subtract=port_4553943c_-port_5a6712aa_;
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_5d300b1c_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_5d300b1c_instance(.GO(GO), 
  .port_5a5faf0f_({subtract[15], subtract[15:1]}), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_5d300b1c_instance_RESULT));
assign RESULT=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_5d300b1c_instance_RESULT;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_5d300b1c_(GO, port_5a5faf0f_, RESULT);
input		GO;
input	[15:0]	port_5a5faf0f_;
output	[15:0]	RESULT;
wire		greaterThan;
wire signed	[15:0]	greaterThan_a_signed;
wire signed	[15:0]	greaterThan_b_signed;
wire		and_u991_u0;
wire		not_u215_u0;
wire		and_u992_u0;
wire		and_u993_u0;
wire	[15:0]	mux_u60;
wire		and_u994_u0;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_5a5faf0f_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign and_u991_u0=GO&not_u215_u0;
assign not_u215_u0=~greaterThan;
assign and_u992_u0=GO&greaterThan;
assign and_u993_u0=and_u992_u0&GO;
assign mux_u60=(and_u994_u0)?port_5a5faf0f_:16'h0;
assign and_u994_u0=and_u991_u0&GO;
assign RESULT=mux_u60;
endmodule



module LL1_L_iunzipFilter2D_midLeftNoConsume2(CLK, RESET, GO, port_056011bc_, port_535b0b03_, port_383828d2_, port_1ffe318b_, RESULT, RESULT_u474, RESULT_u475, RESULT_u476, RESULT_u477, RESULT_u478, RESULT_u479, RESULT_u480, RESULT_u481, RESULT_u482, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_056011bc_;
input	[15:0]	port_535b0b03_;
input		port_383828d2_;
input	[15:0]	port_1ffe318b_;
output		RESULT;
output	[15:0]	RESULT_u474;
output		RESULT_u475;
output	[15:0]	RESULT_u476;
output		RESULT_u477;
output	[31:0]	RESULT_u478;
output	[2:0]	RESULT_u479;
output	[15:0]	RESULT_u480;
output		RESULT_u481;
output	[15:0]	RESULT_u482;
output		DONE;
reg		done_cache_u48=1'h0;
wire		and_u998_u0;
wire		or_u274_u0;
wire		or_u275_u0;
wire		and_u1003_u0;
reg		done_cache_u49_u0=1'h0;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_54b9665a_instance_RESULT;
wire	[15:0]	add;
wire		simplePinWrite;
wire	[15:0]	simplePinWrite_u157;
wire	[15:0]	simplePinWrite_u158;
reg		reg_6503f612_u0=1'h0;
reg	[15:0]	syncEnable_u36=16'h0;
reg		reg_2e9f34be_u0=1'h0;
reg		reg_6503f612_result_delayed_u0=1'h0;
wire		or_u276_u0;
reg		reg_2e9f34be_result_delayed_u0=1'h0;
reg		reg_60857645_u0=1'h0;
always @(posedge CLK or posedge GO or posedge or_u274_u0)
begin
if (or_u274_u0)
done_cache_u48<=1'h0;
else if (GO)
done_cache_u48<=1'h1;
else done_cache_u48<=done_cache_u48;
end
assign and_u998_u0=done_cache_u48&port_383828d2_;
assign or_u274_u0=and_u998_u0|RESET;
assign or_u275_u0=and_u1003_u0|RESET;
assign and_u1003_u0=done_cache_u49_u0&port_383828d2_;
always @(posedge CLK or posedge reg_2e9f34be_u0 or posedge or_u275_u0)
begin
if (or_u275_u0)
done_cache_u49_u0<=1'h0;
else if (reg_2e9f34be_u0)
done_cache_u49_u0<=1'h1;
else done_cache_u49_u0<=done_cache_u49_u0;
end
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_54b9665a_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_54b9665a_instance(.GO(reg_2e9f34be_result_delayed_u0), 
  .port_4a46e936_(port_1ffe318b_), .port_389e3ef6_(syncEnable_u36), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_54b9665a_instance_RESULT));
assign add=port_535b0b03_+16'h1;
assign simplePinWrite=reg_2e9f34be_result_delayed_u0&{1{reg_2e9f34be_result_delayed_u0}};
assign simplePinWrite_u157=16'h1&{16{1'h1}};
assign simplePinWrite_u158=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_54b9665a_instance_RESULT&{16{reg_2e9f34be_result_delayed_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6503f612_u0<=1'h0;
else reg_6503f612_u0<=reg_2e9f34be_result_delayed_u0;
end
always @(posedge CLK)
begin
if (reg_60857645_u0)
syncEnable_u36<=port_1ffe318b_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2e9f34be_u0<=1'h0;
else reg_2e9f34be_u0<=reg_60857645_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6503f612_result_delayed_u0<=1'h0;
else reg_6503f612_result_delayed_u0<=reg_6503f612_u0;
end
assign or_u276_u0=GO|reg_2e9f34be_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2e9f34be_result_delayed_u0<=1'h0;
else reg_2e9f34be_result_delayed_u0<=reg_2e9f34be_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_60857645_u0<=1'h0;
else reg_60857645_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u474=16'h0;
assign RESULT_u475=GO;
assign RESULT_u476=add;
assign RESULT_u477=or_u276_u0;
assign RESULT_u478=32'h0;
assign RESULT_u479=3'h1;
assign RESULT_u480=simplePinWrite_u158;
assign RESULT_u481=simplePinWrite;
assign RESULT_u482=simplePinWrite_u157;
assign DONE=reg_6503f612_result_delayed_u0;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_54b9665a_(GO, port_4a46e936_, port_389e3ef6_, RESULT);
input		GO;
input	[15:0]	port_4a46e936_;
input	[15:0]	port_389e3ef6_;
output	[15:0]	RESULT;
wire	[15:0]	subtract;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_1e6fcbe9_instance_RESULT;
assign subtract=port_389e3ef6_-port_4a46e936_;
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_1e6fcbe9_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_1e6fcbe9_instance(.GO(GO), 
  .port_7305ae3f_({subtract[15], subtract[15:1]}), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_1e6fcbe9_instance_RESULT));
assign RESULT=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_1e6fcbe9_instance_RESULT;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_1e6fcbe9_(GO, port_7305ae3f_, RESULT);
input		GO;
input	[15:0]	port_7305ae3f_;
output	[15:0]	RESULT;
wire		greaterThan;
wire signed	[15:0]	greaterThan_a_signed;
wire signed	[15:0]	greaterThan_b_signed;
wire		and_u1007_u0;
wire		and_u1008_u0;
wire		not_u216_u0;
wire		and_u1009_u0;
wire		and_u1010_u0;
wire	[15:0]	mux_u61;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_7305ae3f_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign and_u1007_u0=GO&not_u216_u0;
assign and_u1008_u0=GO&greaterThan;
assign not_u216_u0=~greaterThan;
assign and_u1009_u0=and_u1007_u0&GO;
assign and_u1010_u0=and_u1008_u0&GO;
assign mux_u61=(and_u1010_u0)?16'h0:port_7305ae3f_;
assign RESULT=mux_u61;
endmodule



module LL1_L_iunzipFilter2D_bottomLeftNoConsume2(CLK, RESET, GO, port_14deb7ac_, port_68ceecfc_, port_3f625033_, port_1c9ca6f6_, RESULT, RESULT_u483, RESULT_u484, RESULT_u485, RESULT_u486, RESULT_u487, RESULT_u488, RESULT_u489, RESULT_u490, RESULT_u491, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_14deb7ac_;
input	[15:0]	port_68ceecfc_;
input		port_3f625033_;
input	[15:0]	port_1c9ca6f6_;
output		RESULT;
output	[15:0]	RESULT_u483;
output		RESULT_u484;
output	[15:0]	RESULT_u485;
output		RESULT_u486;
output	[31:0]	RESULT_u487;
output	[2:0]	RESULT_u488;
output	[15:0]	RESULT_u489;
output	[15:0]	RESULT_u490;
output		RESULT_u491;
output		DONE;
wire		or_u277_u0;
reg		done_cache_u50=1'h0;
wire		and_u1012_u0;
wire		or_u278_u0;
wire		and_u1017_u0;
reg		done_cache_u51_u0=1'h0;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_347f6246_instance_RESULT;
wire	[15:0]	add;
wire	[15:0]	simplePinWrite;
wire	[15:0]	simplePinWrite_u159;
wire		simplePinWrite_u160;
reg		reg_72aa07b2_u0=1'h0;
wire		or_u279_u0;
reg		reg_4e58d7dd_u0=1'h0;
reg	[15:0]	syncEnable_u37=16'h0;
reg		reg_3bcbab60_u0=1'h0;
reg		reg_52bcd111_u0=1'h0;
reg		reg_4e58d7dd_result_delayed_u0=1'h0;
assign or_u277_u0=and_u1012_u0|RESET;
always @(posedge CLK or posedge GO or posedge or_u277_u0)
begin
if (or_u277_u0)
done_cache_u50<=1'h0;
else if (GO)
done_cache_u50<=1'h1;
else done_cache_u50<=done_cache_u50;
end
assign and_u1012_u0=done_cache_u50&port_3f625033_;
assign or_u278_u0=and_u1017_u0|RESET;
assign and_u1017_u0=done_cache_u51_u0&port_3f625033_;
always @(posedge CLK or posedge reg_4e58d7dd_u0 or posedge or_u278_u0)
begin
if (or_u278_u0)
done_cache_u51_u0<=1'h0;
else if (reg_4e58d7dd_u0)
done_cache_u51_u0<=1'h1;
else done_cache_u51_u0<=done_cache_u51_u0;
end
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_347f6246_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_347f6246_instance(.GO(reg_4e58d7dd_result_delayed_u0), 
  .port_62d4d4e4_(port_1c9ca6f6_), .port_585c4360_(syncEnable_u37), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_347f6246_instance_RESULT));
assign add=port_68ceecfc_+16'h1;
assign simplePinWrite=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_347f6246_instance_RESULT&{16{reg_4e58d7dd_result_delayed_u0}};
assign simplePinWrite_u159=16'h1&{16{1'h1}};
assign simplePinWrite_u160=reg_4e58d7dd_result_delayed_u0&{1{reg_4e58d7dd_result_delayed_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_72aa07b2_u0<=1'h0;
else reg_72aa07b2_u0<=reg_52bcd111_u0;
end
assign or_u279_u0=GO|reg_4e58d7dd_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4e58d7dd_u0<=1'h0;
else reg_4e58d7dd_u0<=reg_3bcbab60_u0;
end
always @(posedge CLK)
begin
if (reg_3bcbab60_u0)
syncEnable_u37<=port_1c9ca6f6_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3bcbab60_u0<=1'h0;
else reg_3bcbab60_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_52bcd111_u0<=1'h0;
else reg_52bcd111_u0<=reg_4e58d7dd_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4e58d7dd_result_delayed_u0<=1'h0;
else reg_4e58d7dd_result_delayed_u0<=reg_4e58d7dd_u0;
end
assign RESULT=GO;
assign RESULT_u483=16'h0;
assign RESULT_u484=GO;
assign RESULT_u485=add;
assign RESULT_u486=or_u279_u0;
assign RESULT_u487=32'h0;
assign RESULT_u488=3'h1;
assign RESULT_u489=simplePinWrite;
assign RESULT_u490=simplePinWrite_u159;
assign RESULT_u491=simplePinWrite_u160;
assign DONE=reg_72aa07b2_u0;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_347f6246_(GO, port_62d4d4e4_, port_585c4360_, RESULT);
input		GO;
input	[15:0]	port_62d4d4e4_;
input	[15:0]	port_585c4360_;
output	[15:0]	RESULT;
wire	[15:0]	subtract;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_699d8e81_instance_RESULT;
assign subtract=port_585c4360_-port_62d4d4e4_;
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_699d8e81_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_699d8e81_instance(.GO(GO), 
  .port_1638d6f1_({subtract[15], subtract[15:1]}), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_699d8e81_instance_RESULT));
assign RESULT=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_699d8e81_instance_RESULT;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_699d8e81_(GO, port_1638d6f1_, RESULT);
input		GO;
input	[15:0]	port_1638d6f1_;
output	[15:0]	RESULT;
wire		greaterThan;
wire signed	[15:0]	greaterThan_a_signed;
wire signed	[15:0]	greaterThan_b_signed;
wire		not_u217_u0;
wire		and_u1021_u0;
wire		and_u1022_u0;
wire		and_u1023_u0;
wire	[15:0]	mux_u62;
wire		and_u1024_u0;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_1638d6f1_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign not_u217_u0=~greaterThan;
assign and_u1021_u0=GO&not_u217_u0;
assign and_u1022_u0=GO&greaterThan;
assign and_u1023_u0=and_u1022_u0&GO;
assign mux_u62=(and_u1023_u0)?16'h0:port_1638d6f1_;
assign and_u1024_u0=and_u1021_u0&GO;
assign RESULT=mux_u62;
endmodule



module LL1_L_iunzipFilter2D_topRow(CLK, RESET, GO, port_47a9ee1b_, port_6d5aabbe_, port_1f199a95_, port_2297a1f9_, port_7ad5e7a2_, port_7f824f8f_, port_63075f82_, RESULT, RESULT_u492, RESULT_u493, RESULT_u494, RESULT_u495, RESULT_u496, RESULT_u497, RESULT_u498, RESULT_u499, RESULT_u500, RESULT_u501, RESULT_u502, RESULT_u503, RESULT_u504, RESULT_u505, RESULT_u506, RESULT_u507, RESULT_u508, RESULT_u509, DONE);
input		CLK;
input		RESET;
input		GO;
input	[31:0]	port_47a9ee1b_;
input	[15:0]	port_6d5aabbe_;
input	[15:0]	port_1f199a95_;
input		port_2297a1f9_;
input	[15:0]	port_7ad5e7a2_;
input		port_7f824f8f_;
input	[15:0]	port_63075f82_;
output		RESULT;
output	[31:0]	RESULT_u492;
output		RESULT_u493;
output	[15:0]	RESULT_u494;
output		RESULT_u495;
output	[15:0]	RESULT_u496;
output		RESULT_u497;
output	[15:0]	RESULT_u498;
output		RESULT_u499;
output	[31:0]	RESULT_u500;
output	[2:0]	RESULT_u501;
output		RESULT_u502;
output	[31:0]	RESULT_u503;
output	[15:0]	RESULT_u504;
output	[2:0]	RESULT_u505;
output	[15:0]	RESULT_u506;
output	[15:0]	RESULT_u507;
output		RESULT_u508;
output		RESULT_u509;
output		DONE;
wire		simplePinWrite;
reg		done_cache_u52=1'h0;
wire		and_u1027_u0;
wire		or_u280_u0;
reg		done_cache_u53_u0=1'h0;
wire		and_u1031_u0;
wire		or_u281_u0;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_47251712_instance_RESULT;
wire		or_u282_u0;
wire		and_u1040_u0;
reg		reg_07e6f0d9_u0=1'h0;
wire	[31:0]	add;
wire	[15:0]	add_u13;
wire	[15:0]	add_u14;
wire	[15:0]	simplePinWrite_u161;
wire	[15:0]	simplePinWrite_u162;
wire		simplePinWrite_u163;
reg	[15:0]	syncEnable_u38=16'h0;
reg		reg_4fd7588a_u0=1'h0;
reg		reg_6340fbcf_u0=1'h0;
reg		reg_4fd7588a_result_delayed_u0=1'h0;
reg	[15:0]	syncEnable_u39_u0=16'h0;
wire		or_u283_u0;
reg		reg_05512ebe_u0=1'h0;
reg		reg_1e0feaf9_u0=1'h0;
reg		reg_4fd7588a_result_delayed_result_delayed_u0=1'h0;
assign simplePinWrite=GO&{1{GO}};
always @(posedge CLK or posedge GO or posedge or_u280_u0)
begin
if (or_u280_u0)
done_cache_u52<=1'h0;
else if (GO)
done_cache_u52<=1'h1;
else done_cache_u52<=done_cache_u52;
end
assign and_u1027_u0=done_cache_u52&port_7f824f8f_;
assign or_u280_u0=and_u1027_u0|RESET;
always @(posedge CLK or posedge reg_6340fbcf_u0 or posedge or_u281_u0)
begin
if (or_u281_u0)
done_cache_u53_u0<=1'h0;
else if (reg_6340fbcf_u0)
done_cache_u53_u0<=1'h1;
else done_cache_u53_u0<=done_cache_u53_u0;
end
assign and_u1031_u0=done_cache_u53_u0&port_7f824f8f_;
assign or_u281_u0=and_u1031_u0|RESET;
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_47251712_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_47251712_instance(.GO(reg_4fd7588a_u0), 
  .port_0e6e1d22_(syncEnable_u39_u0), .port_5258c8fa_(port_7ad5e7a2_), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_47251712_instance_RESULT));
assign or_u282_u0=and_u1040_u0|RESET;
assign and_u1040_u0=reg_07e6f0d9_u0&port_7f824f8f_;
always @(posedge CLK or posedge reg_4fd7588a_result_delayed_result_delayed_u0 or posedge or_u282_u0)
begin
if (or_u282_u0)
reg_07e6f0d9_u0<=1'h0;
else if (reg_4fd7588a_result_delayed_result_delayed_u0)
reg_07e6f0d9_u0<=1'h1;
else reg_07e6f0d9_u0<=reg_07e6f0d9_u0;
end
assign add=port_47a9ee1b_+32'h1;
assign add_u13=port_6d5aabbe_+16'h1;
assign add_u14=port_1f199a95_+16'h1;
assign simplePinWrite_u161=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_47251712_instance_RESULT&{16{reg_4fd7588a_u0}};
assign simplePinWrite_u162=16'h1&{16{1'h1}};
assign simplePinWrite_u163=reg_4fd7588a_u0&{1{reg_4fd7588a_u0}};
always @(posedge CLK)
begin
if (GO)
syncEnable_u38<=port_63075f82_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4fd7588a_u0<=1'h0;
else reg_4fd7588a_u0<=reg_6340fbcf_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6340fbcf_u0<=1'h0;
else reg_6340fbcf_u0<=reg_1e0feaf9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4fd7588a_result_delayed_u0<=1'h0;
else reg_4fd7588a_result_delayed_u0<=reg_4fd7588a_u0;
end
always @(posedge CLK)
begin
if (reg_1e0feaf9_u0)
syncEnable_u39_u0<=port_7ad5e7a2_;
end
assign or_u283_u0=GO|reg_6340fbcf_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_05512ebe_u0<=1'h0;
else reg_05512ebe_u0<=reg_4fd7588a_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1e0feaf9_u0<=1'h0;
else reg_1e0feaf9_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4fd7588a_result_delayed_result_delayed_u0<=1'h0;
else reg_4fd7588a_result_delayed_result_delayed_u0<=reg_4fd7588a_result_delayed_u0;
end
assign RESULT=GO;
assign RESULT_u492=add;
assign RESULT_u493=GO;
assign RESULT_u494=16'h0;
assign RESULT_u495=GO;
assign RESULT_u496=add_u13;
assign RESULT_u497=GO;
assign RESULT_u498=add_u14;
assign RESULT_u499=or_u283_u0;
assign RESULT_u500=32'h0;
assign RESULT_u501=3'h1;
assign RESULT_u502=reg_4fd7588a_result_delayed_result_delayed_u0;
assign RESULT_u503=32'h0;
assign RESULT_u504=syncEnable_u38;
assign RESULT_u505=3'h1;
assign RESULT_u506=simplePinWrite_u161;
assign RESULT_u507=simplePinWrite_u162;
assign RESULT_u508=simplePinWrite;
assign RESULT_u509=simplePinWrite_u163;
assign DONE=reg_05512ebe_u0;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_47251712_(GO, port_0e6e1d22_, port_5258c8fa_, RESULT);
input		GO;
input	[15:0]	port_0e6e1d22_;
input	[15:0]	port_5258c8fa_;
output	[15:0]	RESULT;
wire	[16:0]	add;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_1fa615f7_instance_RESULT;
assign add={port_0e6e1d22_[15], port_0e6e1d22_}+{port_5258c8fa_[15], port_5258c8fa_};
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_1fa615f7_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_1fa615f7_instance(.GO(GO), 
  .port_3626a115_({add[16], add[16:2]}), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_1fa615f7_instance_RESULT));
assign RESULT=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_1fa615f7_instance_RESULT;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_1fa615f7_(GO, port_3626a115_, RESULT);
input		GO;
input	[15:0]	port_3626a115_;
output	[15:0]	RESULT;
wire signed	[15:0]	greaterThan_b_signed;
wire signed	[15:0]	greaterThan_a_signed;
wire		greaterThan;
wire		and_u1035_u0;
wire		and_u1036_u0;
wire		not_u218_u0;
wire	[15:0]	mux_u63;
wire		and_u1037_u0;
wire		and_u1038_u0;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_3626a115_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign and_u1035_u0=GO&greaterThan;
assign and_u1036_u0=GO&not_u218_u0;
assign not_u218_u0=~greaterThan;
assign mux_u63=(and_u1038_u0)?port_3626a115_:16'h0;
assign and_u1037_u0=and_u1035_u0&GO;
assign and_u1038_u0=and_u1036_u0&GO;
assign RESULT=mux_u63;
endmodule



module LL1_L_iunzipFilter2D_endianswapper_33a44bd8_(endianswapper_33a44bd8_in, endianswapper_33a44bd8_out);
input	[15:0]	endianswapper_33a44bd8_in;
output	[15:0]	endianswapper_33a44bd8_out;
assign endianswapper_33a44bd8_out=endianswapper_33a44bd8_in;
endmodule



module LL1_L_iunzipFilter2D_endianswapper_26e2d6fe_(endianswapper_26e2d6fe_in, endianswapper_26e2d6fe_out);
input	[15:0]	endianswapper_26e2d6fe_in;
output	[15:0]	endianswapper_26e2d6fe_out;
assign endianswapper_26e2d6fe_out=endianswapper_26e2d6fe_in;
endmodule



module LL1_L_iunzipFilter2D_stateVar_populatePtr(bus_4bd01fea_, bus_5e5c669f_, bus_5000423d_, bus_2631ddf5_, bus_2160680b_, bus_338c8ca8_, bus_3ae80db9_);
input		bus_4bd01fea_;
input		bus_5e5c669f_;
input		bus_5000423d_;
input	[15:0]	bus_2631ddf5_;
input		bus_2160680b_;
input	[15:0]	bus_338c8ca8_;
output	[15:0]	bus_3ae80db9_;
wire	[15:0]	mux_7765a436_u0;
reg	[15:0]	stateVar_populatePtr_u1=16'h0;
wire		or_58ddc804_u0;
wire	[15:0]	endianswapper_33a44bd8_out;
wire	[15:0]	endianswapper_26e2d6fe_out;
assign mux_7765a436_u0=(bus_5000423d_)?bus_2631ddf5_:16'h0;
always @(posedge bus_4bd01fea_ or posedge bus_5e5c669f_)
begin
if (bus_5e5c669f_)
stateVar_populatePtr_u1<=16'h0;
else if (or_58ddc804_u0)
stateVar_populatePtr_u1<=endianswapper_33a44bd8_out;
end
assign bus_3ae80db9_=endianswapper_26e2d6fe_out;
assign or_58ddc804_u0=bus_5000423d_|bus_2160680b_;
LL1_L_iunzipFilter2D_endianswapper_33a44bd8_ LL1_L_iunzipFilter2D_endianswapper_33a44bd8__1(.endianswapper_33a44bd8_in(mux_7765a436_u0), 
  .endianswapper_33a44bd8_out(endianswapper_33a44bd8_out));
LL1_L_iunzipFilter2D_endianswapper_26e2d6fe_ LL1_L_iunzipFilter2D_endianswapper_26e2d6fe__1(.endianswapper_26e2d6fe_in(stateVar_populatePtr_u1), 
  .endianswapper_26e2d6fe_out(endianswapper_26e2d6fe_out));
endmodule



module LL1_L_iunzipFilter2D_midRight1(CLK, RESET, GO, port_5255d759_, port_14c39ecd_, port_282e491b_, port_4c76bba0_, port_631edf34_, port_2c10671c_, port_07cc4909_, RESULT, RESULT_u510, RESULT_u511, RESULT_u512, RESULT_u513, RESULT_u514, RESULT_u515, RESULT_u516, RESULT_u517, RESULT_u518, RESULT_u519, RESULT_u520, RESULT_u521, RESULT_u522, RESULT_u523, RESULT_u524, RESULT_u525, RESULT_u526, RESULT_u527, RESULT_u528, RESULT_u529, DONE);
input		CLK;
input		RESET;
input		GO;
input	[31:0]	port_5255d759_;
input	[15:0]	port_14c39ecd_;
input		port_282e491b_;
input		port_4c76bba0_;
input	[15:0]	port_631edf34_;
input		port_2c10671c_;
input	[15:0]	port_07cc4909_;
output		RESULT;
output	[15:0]	RESULT_u510;
output		RESULT_u511;
output	[31:0]	RESULT_u512;
output		RESULT_u513;
output	[15:0]	RESULT_u514;
output		RESULT_u515;
output	[15:0]	RESULT_u516;
output		RESULT_u517;
output		RESULT_u518;
output		RESULT_u519;
output	[31:0]	RESULT_u520;
output	[2:0]	RESULT_u521;
output		RESULT_u522;
output	[31:0]	RESULT_u523;
output	[15:0]	RESULT_u524;
output	[2:0]	RESULT_u525;
output	[15:0]	RESULT_u526;
output	[15:0]	RESULT_u527;
output		RESULT_u528;
output		RESULT_u529;
output		DONE;
wire		simplePinWrite;
reg		done_cache_u54=1'h0;
wire		and_u1043_u0;
wire		or_u284_u0;
reg		done_cache_u55_u0=1'h0;
wire		or_u285_u0;
wire		and_u1048_u0;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_39faca6a_instance_RESULT;
wire		and_u1057_u0;
reg		reg_70d2a446_u0=1'h0;
wire		or_u286_u0;
wire	[31:0]	add;
wire	[15:0]	add_u15;
wire		not_u220;
wire	[15:0]	simplePinWrite_u164;
wire		simplePinWrite_u165;
wire	[15:0]	simplePinWrite_u166;
reg		reg_5a9aa882_u0=1'h0;
reg		reg_145a3242_u0=1'h0;
reg		reg_354d1b6c_u0=1'h0;
reg		reg_145a3242_result_delayed_u0=1'h0;
reg	[15:0]	syncEnable_u40=16'h0;
reg	[15:0]	syncEnable_u41_u0=16'h0;
reg		reg_5a9aa882_result_delayed_u0=1'h0;
wire		or_u287_u0;
reg		reg_1b3d28e6_u0=1'h0;
assign simplePinWrite=GO&{1{GO}};
always @(posedge CLK or posedge GO or posedge or_u284_u0)
begin
if (or_u284_u0)
done_cache_u54<=1'h0;
else if (GO)
done_cache_u54<=1'h1;
else done_cache_u54<=done_cache_u54;
end
assign and_u1043_u0=done_cache_u54&port_2c10671c_;
assign or_u284_u0=and_u1043_u0|RESET;
always @(posedge CLK or posedge reg_5a9aa882_u0 or posedge or_u285_u0)
begin
if (or_u285_u0)
done_cache_u55_u0<=1'h0;
else if (reg_5a9aa882_u0)
done_cache_u55_u0<=1'h1;
else done_cache_u55_u0<=done_cache_u55_u0;
end
assign or_u285_u0=and_u1048_u0|RESET;
assign and_u1048_u0=done_cache_u55_u0&port_2c10671c_;
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_39faca6a_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_39faca6a_instance(.GO(reg_5a9aa882_result_delayed_u0), 
  .port_09ce286e_(syncEnable_u40), .port_0e1040f8_(port_631edf34_), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_39faca6a_instance_RESULT));
assign and_u1057_u0=reg_70d2a446_u0&port_2c10671c_;
always @(posedge CLK or posedge reg_145a3242_u0 or posedge or_u286_u0)
begin
if (or_u286_u0)
reg_70d2a446_u0<=1'h0;
else if (reg_145a3242_u0)
reg_70d2a446_u0<=1'h1;
else reg_70d2a446_u0<=reg_70d2a446_u0;
end
assign or_u286_u0=and_u1057_u0|RESET;
assign add=port_5255d759_+32'h1;
assign add_u15=port_14c39ecd_+16'h1;
assign not_u220=!port_282e491b_;
assign simplePinWrite_u164=16'h1&{16{1'h1}};
assign simplePinWrite_u165=reg_5a9aa882_result_delayed_u0&{1{reg_5a9aa882_result_delayed_u0}};
assign simplePinWrite_u166=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_39faca6a_instance_RESULT&{16{reg_5a9aa882_result_delayed_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5a9aa882_u0<=1'h0;
else reg_5a9aa882_u0<=reg_1b3d28e6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_145a3242_u0<=1'h0;
else reg_145a3242_u0<=reg_354d1b6c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_354d1b6c_u0<=1'h0;
else reg_354d1b6c_u0<=reg_5a9aa882_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_145a3242_result_delayed_u0<=1'h0;
else reg_145a3242_result_delayed_u0<=reg_145a3242_u0;
end
always @(posedge CLK)
begin
if (reg_1b3d28e6_u0)
syncEnable_u40<=port_631edf34_;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u41_u0<=port_07cc4909_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5a9aa882_result_delayed_u0<=1'h0;
else reg_5a9aa882_result_delayed_u0<=reg_5a9aa882_u0;
end
assign or_u287_u0=GO|reg_5a9aa882_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1b3d28e6_u0<=1'h0;
else reg_1b3d28e6_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u510=16'h0;
assign RESULT_u511=GO;
assign RESULT_u512=add;
assign RESULT_u513=GO;
assign RESULT_u514=add_u15;
assign RESULT_u515=GO;
assign RESULT_u516=16'h0;
assign RESULT_u517=GO;
assign RESULT_u518=not_u220;
assign RESULT_u519=or_u287_u0;
assign RESULT_u520=32'h0;
assign RESULT_u521=3'h1;
assign RESULT_u522=reg_145a3242_u0;
assign RESULT_u523=32'h0;
assign RESULT_u524=syncEnable_u41_u0;
assign RESULT_u525=3'h1;
assign RESULT_u526=simplePinWrite_u166;
assign RESULT_u527=simplePinWrite_u164;
assign RESULT_u528=simplePinWrite;
assign RESULT_u529=simplePinWrite_u165;
assign DONE=reg_145a3242_result_delayed_u0;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_39faca6a_(GO, port_09ce286e_, port_0e1040f8_, RESULT);
input		GO;
input	[15:0]	port_09ce286e_;
input	[15:0]	port_0e1040f8_;
output	[15:0]	RESULT;
wire	[16:0]	add;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_529aa0aa_instance_RESULT;
assign add={port_09ce286e_[15], port_09ce286e_}+{port_0e1040f8_[15], port_0e1040f8_};
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_529aa0aa_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_529aa0aa_instance(.GO(GO), 
  .port_4a4d51aa_({add[16], add[16:2]}), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_529aa0aa_instance_RESULT));
assign RESULT=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_529aa0aa_instance_RESULT;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_529aa0aa_(GO, port_4a4d51aa_, RESULT);
input		GO;
input	[15:0]	port_4a4d51aa_;
output	[15:0]	RESULT;
wire signed	[15:0]	greaterThan_a_signed;
wire signed	[15:0]	greaterThan_b_signed;
wire		greaterThan;
wire		not_u219_u0;
wire		and_u1052_u0;
wire		and_u1053_u0;
wire		and_u1054_u0;
wire		and_u1055_u0;
wire	[15:0]	mux_u64;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_4a4d51aa_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign not_u219_u0=~greaterThan;
assign and_u1052_u0=GO&greaterThan;
assign and_u1053_u0=GO&not_u219_u0;
assign and_u1054_u0=and_u1053_u0&GO;
assign and_u1055_u0=and_u1052_u0&GO;
assign mux_u64=(and_u1055_u0)?16'h0:port_4a4d51aa_;
assign RESULT=mux_u64;
endmodule



module LL1_L_iunzipFilter2D_stateVar_isEven(bus_1f3489ff_, bus_4d0fbe00_, bus_7316061a_, bus_78994a42_, bus_52631b34_, bus_1823e66f_, bus_743d02cc_, bus_0a184a25_, bus_40103492_, bus_7b46d837_, bus_5dc6e0f1_, bus_1c6f5c87_, bus_75eeb741_, bus_6f55ec5d_, bus_581ab06d_, bus_51887cdb_, bus_6b52f69a_);
input		bus_1f3489ff_;
input		bus_4d0fbe00_;
input		bus_7316061a_;
input		bus_78994a42_;
input		bus_52631b34_;
input		bus_1823e66f_;
input		bus_743d02cc_;
input		bus_0a184a25_;
input		bus_40103492_;
input		bus_7b46d837_;
input		bus_5dc6e0f1_;
input		bus_1c6f5c87_;
input		bus_75eeb741_;
input		bus_6f55ec5d_;
input		bus_581ab06d_;
input		bus_51887cdb_;
output		bus_6b52f69a_;
wire		mux_4262b723_u0;
reg		stateVar_isEven_u1=1'h1;
wire		or_25632e9a_u0;
assign mux_4262b723_u0=({1{bus_7316061a_}}&bus_78994a42_)|({1{bus_52631b34_}}&bus_1823e66f_)|({1{bus_743d02cc_}}&bus_0a184a25_)|({1{bus_40103492_}}&bus_7b46d837_)|({1{bus_5dc6e0f1_}}&bus_1c6f5c87_)|({1{bus_75eeb741_}}&bus_6f55ec5d_)|({1{bus_581ab06d_}}&bus_51887cdb_);
always @(posedge bus_1f3489ff_ or posedge bus_4d0fbe00_)
begin
if (bus_4d0fbe00_)
stateVar_isEven_u1<=1'h1;
else if (or_25632e9a_u0)
stateVar_isEven_u1<=mux_4262b723_u0;
end
assign or_25632e9a_u0=bus_7316061a_|bus_52631b34_|bus_743d02cc_|bus_40103492_|bus_5dc6e0f1_|bus_75eeb741_|bus_581ab06d_;
assign bus_6b52f69a_=stateVar_isEven_u1;
endmodule



module LL1_L_iunzipFilter2D_midRight2(CLK, RESET, GO, port_7204953c_, port_1cd54e3f_, port_2166078e_, port_38854079_, port_1fe65f07_, port_2a04576f_, port_6e163b29_, RESULT, RESULT_u530, RESULT_u531, RESULT_u532, RESULT_u533, RESULT_u534, RESULT_u535, RESULT_u536, RESULT_u537, RESULT_u538, RESULT_u539, RESULT_u540, RESULT_u541, RESULT_u542, RESULT_u543, RESULT_u544, RESULT_u545, RESULT_u546, RESULT_u547, RESULT_u548, RESULT_u549, DONE);
input		CLK;
input		RESET;
input		GO;
input	[31:0]	port_7204953c_;
input	[15:0]	port_1cd54e3f_;
input		port_2166078e_;
input		port_38854079_;
input	[15:0]	port_1fe65f07_;
input		port_2a04576f_;
input	[15:0]	port_6e163b29_;
output		RESULT;
output	[15:0]	RESULT_u530;
output		RESULT_u531;
output	[31:0]	RESULT_u532;
output		RESULT_u533;
output	[15:0]	RESULT_u534;
output		RESULT_u535;
output	[15:0]	RESULT_u536;
output		RESULT_u537;
output		RESULT_u538;
output		RESULT_u539;
output	[31:0]	RESULT_u540;
output	[2:0]	RESULT_u541;
output		RESULT_u542;
output	[31:0]	RESULT_u543;
output	[15:0]	RESULT_u544;
output	[2:0]	RESULT_u545;
output	[15:0]	RESULT_u546;
output		RESULT_u547;
output		RESULT_u548;
output	[15:0]	RESULT_u549;
output		DONE;
wire		simplePinWrite;
wire		and_u1060_u0;
wire		or_u288_u0;
reg		done_cache_u56=1'h0;
wire		or_u289_u0;
reg		done_cache_u57_u0=1'h0;
wire		and_u1065_u0;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_16f9a1af_instance_RESULT;
reg		reg_5bcbf79f_u0=1'h0;
wire		or_u290_u0;
wire		and_u1074_u0;
wire	[31:0]	add;
wire	[15:0]	add_u16;
wire		not_u222;
wire	[15:0]	simplePinWrite_u167;
wire		simplePinWrite_u168;
wire	[15:0]	simplePinWrite_u169;
reg		reg_23df0fab_u0=1'h0;
reg		reg_5c3e96b6_u0=1'h0;
reg		reg_73247d86_u0=1'h0;
wire		or_u291_u0;
reg		reg_632073c9_u0=1'h0;
reg	[15:0]	syncEnable_u42=16'h0;
reg		reg_1edea7ae_u0=1'h0;
reg		reg_23df0fab_result_delayed_u0=1'h0;
reg	[15:0]	syncEnable_u43_u0=16'h0;
assign simplePinWrite=GO&{1{GO}};
assign and_u1060_u0=done_cache_u56&port_2a04576f_;
assign or_u288_u0=and_u1060_u0|RESET;
always @(posedge CLK or posedge GO or posedge or_u288_u0)
begin
if (or_u288_u0)
done_cache_u56<=1'h0;
else if (GO)
done_cache_u56<=1'h1;
else done_cache_u56<=done_cache_u56;
end
assign or_u289_u0=and_u1065_u0|RESET;
always @(posedge CLK or posedge reg_73247d86_u0 or posedge or_u289_u0)
begin
if (or_u289_u0)
done_cache_u57_u0<=1'h0;
else if (reg_73247d86_u0)
done_cache_u57_u0<=1'h1;
else done_cache_u57_u0<=done_cache_u57_u0;
end
assign and_u1065_u0=done_cache_u57_u0&port_2a04576f_;
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_16f9a1af_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_16f9a1af_instance(.GO(reg_5c3e96b6_u0), 
  .port_26c781b2_(port_1fe65f07_), .port_17d44117_(syncEnable_u43_u0), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_16f9a1af_instance_RESULT));
always @(posedge CLK or posedge reg_23df0fab_result_delayed_u0 or posedge or_u290_u0)
begin
if (or_u290_u0)
reg_5bcbf79f_u0<=1'h0;
else if (reg_23df0fab_result_delayed_u0)
reg_5bcbf79f_u0<=1'h1;
else reg_5bcbf79f_u0<=reg_5bcbf79f_u0;
end
assign or_u290_u0=and_u1074_u0|RESET;
assign and_u1074_u0=reg_5bcbf79f_u0&port_2a04576f_;
assign add=port_7204953c_+32'h1;
assign add_u16=port_1cd54e3f_+16'h1;
assign not_u222=!port_2166078e_;
assign simplePinWrite_u167=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_16f9a1af_instance_RESULT&{16{reg_5c3e96b6_u0}};
assign simplePinWrite_u168=reg_5c3e96b6_u0&{1{reg_5c3e96b6_u0}};
assign simplePinWrite_u169=16'h1&{16{1'h1}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_23df0fab_u0<=1'h0;
else reg_23df0fab_u0<=reg_5c3e96b6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5c3e96b6_u0<=1'h0;
else reg_5c3e96b6_u0<=reg_73247d86_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_73247d86_u0<=1'h0;
else reg_73247d86_u0<=reg_1edea7ae_u0;
end
assign or_u291_u0=GO|reg_73247d86_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_632073c9_u0<=1'h0;
else reg_632073c9_u0<=reg_23df0fab_result_delayed_u0;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u42<=port_6e163b29_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1edea7ae_u0<=1'h0;
else reg_1edea7ae_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_23df0fab_result_delayed_u0<=1'h0;
else reg_23df0fab_result_delayed_u0<=reg_23df0fab_u0;
end
always @(posedge CLK)
begin
if (reg_1edea7ae_u0)
syncEnable_u43_u0<=port_1fe65f07_;
end
assign RESULT=GO;
assign RESULT_u530=16'h0;
assign RESULT_u531=GO;
assign RESULT_u532=add;
assign RESULT_u533=GO;
assign RESULT_u534=add_u16;
assign RESULT_u535=GO;
assign RESULT_u536=16'h0;
assign RESULT_u537=GO;
assign RESULT_u538=not_u222;
assign RESULT_u539=or_u291_u0;
assign RESULT_u540=32'h0;
assign RESULT_u541=3'h1;
assign RESULT_u542=reg_23df0fab_result_delayed_u0;
assign RESULT_u543=32'h0;
assign RESULT_u544=syncEnable_u42;
assign RESULT_u545=3'h1;
assign RESULT_u546=simplePinWrite_u167;
assign RESULT_u547=simplePinWrite;
assign RESULT_u548=simplePinWrite_u168;
assign RESULT_u549=simplePinWrite_u169;
assign DONE=reg_632073c9_u0;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_16f9a1af_(GO, port_26c781b2_, port_17d44117_, RESULT);
input		GO;
input	[15:0]	port_26c781b2_;
input	[15:0]	port_17d44117_;
output	[15:0]	RESULT;
wire	[15:0]	subtract;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_78e4beec_instance_RESULT;
assign subtract=port_17d44117_-port_26c781b2_;
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_78e4beec_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_78e4beec_instance(.GO(GO), 
  .port_440f8a09_({subtract[15], subtract[15:1]}), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_78e4beec_instance_RESULT));
assign RESULT=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_78e4beec_instance_RESULT;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_78e4beec_(GO, port_440f8a09_, RESULT);
input		GO;
input	[15:0]	port_440f8a09_;
output	[15:0]	RESULT;
wire		greaterThan;
wire signed	[15:0]	greaterThan_a_signed;
wire signed	[15:0]	greaterThan_b_signed;
wire		not_u221_u0;
wire		and_u1069_u0;
wire		and_u1070_u0;
wire		and_u1071_u0;
wire		and_u1072_u0;
wire	[15:0]	mux_u65;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_440f8a09_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign not_u221_u0=~greaterThan;
assign and_u1069_u0=GO&greaterThan;
assign and_u1070_u0=GO&not_u221_u0;
assign and_u1071_u0=and_u1070_u0&GO;
assign and_u1072_u0=and_u1069_u0&GO;
assign mux_u65=(and_u1072_u0)?16'h0:port_440f8a09_;
assign RESULT=mux_u65;
endmodule



module LL1_L_iunzipFilter2D_midLeft1(CLK, RESET, GO, port_250e58ba_, port_6197b3d4_, port_43ef7bd5_, port_36b60040_, port_78b91e36_, port_5a4c347c_, port_616f0feb_, RESULT, RESULT_u550, RESULT_u551, RESULT_u552, RESULT_u553, RESULT_u554, RESULT_u555, RESULT_u556, RESULT_u557, RESULT_u558, RESULT_u559, RESULT_u560, RESULT_u561, RESULT_u562, RESULT_u563, RESULT_u564, RESULT_u565, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_250e58ba_;
input	[31:0]	port_6197b3d4_;
input	[15:0]	port_43ef7bd5_;
input		port_36b60040_;
input	[15:0]	port_78b91e36_;
input		port_5a4c347c_;
input	[15:0]	port_616f0feb_;
output		RESULT;
output	[15:0]	RESULT_u550;
output		RESULT_u551;
output	[31:0]	RESULT_u552;
output		RESULT_u553;
output	[15:0]	RESULT_u554;
output		RESULT_u555;
output	[31:0]	RESULT_u556;
output	[2:0]	RESULT_u557;
output		RESULT_u558;
output	[31:0]	RESULT_u559;
output	[15:0]	RESULT_u560;
output	[2:0]	RESULT_u561;
output	[15:0]	RESULT_u562;
output	[15:0]	RESULT_u563;
output		RESULT_u564;
output		RESULT_u565;
output		DONE;
wire		simplePinWrite;
wire		or_u292_u0;
reg		done_cache_u58=1'h0;
wire		and_u1076_u0;
wire		or_u293_u0;
reg		done_cache_u59_u0=1'h0;
wire		and_u1081_u0;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_57113ac8_instance_RESULT;
wire		or_u294_u0;
wire		and_u1090_u0;
reg		reg_388bdee4_u0=1'h0;
wire	[31:0]	add;
wire	[15:0]	add_u17;
wire	[15:0]	simplePinWrite_u170;
wire	[15:0]	simplePinWrite_u171;
wire		simplePinWrite_u172;
reg		reg_3139452e_u0=1'h0;
reg		reg_3d3b006d_u0=1'h0;
reg	[15:0]	syncEnable_u44=16'h0;
reg		reg_71109e8c_u0=1'h0;
reg		reg_67a8b519_u0=1'h0;
reg	[15:0]	syncEnable_u45_u0=16'h0;
reg		reg_71109e8c_result_delayed_u0=1'h0;
reg		reg_3139452e_result_delayed_u0=1'h0;
wire		or_u295_u0;
assign simplePinWrite=GO&{1{GO}};
assign or_u292_u0=and_u1076_u0|RESET;
always @(posedge CLK or posedge GO or posedge or_u292_u0)
begin
if (or_u292_u0)
done_cache_u58<=1'h0;
else if (GO)
done_cache_u58<=1'h1;
else done_cache_u58<=done_cache_u58;
end
assign and_u1076_u0=done_cache_u58&port_5a4c347c_;
assign or_u293_u0=and_u1081_u0|RESET;
always @(posedge CLK or posedge reg_71109e8c_result_delayed_u0 or posedge or_u293_u0)
begin
if (or_u293_u0)
done_cache_u59_u0<=1'h0;
else if (reg_71109e8c_result_delayed_u0)
done_cache_u59_u0<=1'h1;
else done_cache_u59_u0<=done_cache_u59_u0;
end
assign and_u1081_u0=done_cache_u59_u0&port_5a4c347c_;
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_57113ac8_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_57113ac8_instance(.GO(reg_67a8b519_u0), 
  .port_674873a6_(syncEnable_u45_u0), .port_11d7bd51_(port_78b91e36_), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_57113ac8_instance_RESULT));
assign or_u294_u0=and_u1090_u0|RESET;
assign and_u1090_u0=reg_388bdee4_u0&port_5a4c347c_;
always @(posedge CLK or posedge reg_3139452e_result_delayed_u0 or posedge or_u294_u0)
begin
if (or_u294_u0)
reg_388bdee4_u0<=1'h0;
else if (reg_3139452e_result_delayed_u0)
reg_388bdee4_u0<=1'h1;
else reg_388bdee4_u0<=reg_388bdee4_u0;
end
assign add=port_6197b3d4_+32'h1;
assign add_u17=port_43ef7bd5_+16'h1;
assign simplePinWrite_u170=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_57113ac8_instance_RESULT&{16{reg_67a8b519_u0}};
assign simplePinWrite_u171=16'h1&{16{1'h1}};
assign simplePinWrite_u172=reg_67a8b519_u0&{1{reg_67a8b519_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3139452e_u0<=1'h0;
else reg_3139452e_u0<=reg_67a8b519_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3d3b006d_u0<=1'h0;
else reg_3d3b006d_u0<=reg_3139452e_result_delayed_u0;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u44<=port_616f0feb_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_71109e8c_u0<=1'h0;
else reg_71109e8c_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_67a8b519_u0<=1'h0;
else reg_67a8b519_u0<=reg_71109e8c_result_delayed_u0;
end
always @(posedge CLK)
begin
if (reg_71109e8c_u0)
syncEnable_u45_u0<=port_78b91e36_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_71109e8c_result_delayed_u0<=1'h0;
else reg_71109e8c_result_delayed_u0<=reg_71109e8c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3139452e_result_delayed_u0<=1'h0;
else reg_3139452e_result_delayed_u0<=reg_3139452e_u0;
end
assign or_u295_u0=GO|reg_71109e8c_result_delayed_u0;
assign RESULT=GO;
assign RESULT_u550=16'h0;
assign RESULT_u551=GO;
assign RESULT_u552=add;
assign RESULT_u553=GO;
assign RESULT_u554=add_u17;
assign RESULT_u555=or_u295_u0;
assign RESULT_u556=32'h0;
assign RESULT_u557=3'h1;
assign RESULT_u558=reg_3139452e_result_delayed_u0;
assign RESULT_u559=32'h0;
assign RESULT_u560=syncEnable_u44;
assign RESULT_u561=3'h1;
assign RESULT_u562=simplePinWrite_u170;
assign RESULT_u563=simplePinWrite_u171;
assign RESULT_u564=simplePinWrite;
assign RESULT_u565=simplePinWrite_u172;
assign DONE=reg_3d3b006d_u0;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_57113ac8_(GO, port_674873a6_, port_11d7bd51_, RESULT);
input		GO;
input	[15:0]	port_674873a6_;
input	[15:0]	port_11d7bd51_;
output	[15:0]	RESULT;
wire	[16:0]	add;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_2f5c4a4b_instance_RESULT;
assign add={port_674873a6_[15], port_674873a6_}+{port_11d7bd51_[15], port_11d7bd51_};
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_2f5c4a4b_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_2f5c4a4b_instance(.GO(GO), 
  .port_32cb0240_({add[16], add[16:2]}), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_2f5c4a4b_instance_RESULT));
assign RESULT=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_2f5c4a4b_instance_RESULT;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_2f5c4a4b_(GO, port_32cb0240_, RESULT);
input		GO;
input	[15:0]	port_32cb0240_;
output	[15:0]	RESULT;
wire		greaterThan;
wire signed	[15:0]	greaterThan_a_signed;
wire signed	[15:0]	greaterThan_b_signed;
wire		not_u223_u0;
wire		and_u1085_u0;
wire		and_u1086_u0;
wire	[15:0]	mux_u66;
wire		and_u1087_u0;
wire		and_u1088_u0;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_32cb0240_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign not_u223_u0=~greaterThan;
assign and_u1085_u0=GO&greaterThan;
assign and_u1086_u0=GO&not_u223_u0;
assign mux_u66=(and_u1088_u0)?16'h0:port_32cb0240_;
assign and_u1087_u0=and_u1086_u0&GO;
assign and_u1088_u0=and_u1085_u0&GO;
assign RESULT=mux_u66;
endmodule



module LL1_L_iunzipFilter2D_endianswapper_712f4033_(endianswapper_712f4033_in, endianswapper_712f4033_out);
input	[15:0]	endianswapper_712f4033_in;
output	[15:0]	endianswapper_712f4033_out;
assign endianswapper_712f4033_out=16'h0;
endmodule



module LL1_L_iunzipFilter2D_endianswapper_42c2e6ef_(endianswapper_42c2e6ef_in, endianswapper_42c2e6ef_out);
input	[15:0]	endianswapper_42c2e6ef_in;
output	[15:0]	endianswapper_42c2e6ef_out;
assign endianswapper_42c2e6ef_out=16'h0;
endmodule



module LL1_L_iunzipFilter2D_stateVar_idx(bus_62860c78_, bus_744fb394_, bus_55af70f4_, bus_0ec28381_, bus_7a64655b_, bus_25e2c4f7_, bus_3c68edfe_, bus_04039d41_, bus_6208d411_, bus_6483ddbc_, bus_7f2a89e4_, bus_6cd25c20_, bus_2fe413a1_, bus_77a210b0_, bus_2ad73ea4_, bus_3f7de95e_, bus_0387bc2f_, bus_61448fc8_, bus_7b1a01ba_, bus_12d790ff_, bus_69a6a217_, bus_539c4f12_, bus_1e9c9e19_, bus_4104bb04_, bus_48c5d111_, bus_50263840_, bus_1b1b4f63_, bus_3d8d462c_, bus_03c74654_, bus_4c32e0b1_, bus_0420cb9d_, bus_0f0be065_, bus_563eebef_, bus_6fc1dd73_, bus_1fe6e51c_, bus_09922e92_, bus_2fd9f75a_, bus_153933ae_, bus_0b1e2e3f_, bus_61c6e306_, bus_79ca6720_);
input		bus_62860c78_;
input		bus_744fb394_;
input		bus_55af70f4_;
input	[15:0]	bus_0ec28381_;
input		bus_7a64655b_;
input	[15:0]	bus_25e2c4f7_;
input		bus_3c68edfe_;
input	[15:0]	bus_04039d41_;
input		bus_6208d411_;
input	[15:0]	bus_6483ddbc_;
input		bus_7f2a89e4_;
input	[15:0]	bus_6cd25c20_;
input		bus_2fe413a1_;
input	[15:0]	bus_77a210b0_;
input		bus_2ad73ea4_;
input	[15:0]	bus_3f7de95e_;
input		bus_0387bc2f_;
input	[15:0]	bus_61448fc8_;
input		bus_7b1a01ba_;
input	[15:0]	bus_12d790ff_;
input		bus_69a6a217_;
input	[15:0]	bus_539c4f12_;
input		bus_1e9c9e19_;
input	[15:0]	bus_4104bb04_;
input		bus_48c5d111_;
input	[15:0]	bus_50263840_;
input		bus_1b1b4f63_;
input	[15:0]	bus_3d8d462c_;
input		bus_03c74654_;
input	[15:0]	bus_4c32e0b1_;
input		bus_0420cb9d_;
input	[15:0]	bus_0f0be065_;
input		bus_563eebef_;
input	[15:0]	bus_6fc1dd73_;
input		bus_1fe6e51c_;
input	[15:0]	bus_09922e92_;
input		bus_2fd9f75a_;
input	[15:0]	bus_153933ae_;
input		bus_0b1e2e3f_;
input	[15:0]	bus_61c6e306_;
output	[15:0]	bus_79ca6720_;
wire		or_5a65bb52_u0;
wire	[15:0]	endianswapper_712f4033_out;
wire	[15:0]	endianswapper_42c2e6ef_out;
assign or_5a65bb52_u0=bus_55af70f4_|bus_7a64655b_|bus_3c68edfe_|bus_6208d411_|bus_7f2a89e4_|bus_2fe413a1_|bus_2ad73ea4_|bus_0387bc2f_|bus_7b1a01ba_|bus_69a6a217_|bus_1e9c9e19_|bus_48c5d111_|bus_1b1b4f63_|bus_03c74654_|bus_0420cb9d_|bus_563eebef_|bus_1fe6e51c_|bus_2fd9f75a_|bus_0b1e2e3f_;
assign bus_79ca6720_=16'h0;
LL1_L_iunzipFilter2D_endianswapper_712f4033_ LL1_L_iunzipFilter2D_endianswapper_712f4033__1(.endianswapper_712f4033_in(16'h0), 
  .endianswapper_712f4033_out(endianswapper_712f4033_out));
LL1_L_iunzipFilter2D_endianswapper_42c2e6ef_ LL1_L_iunzipFilter2D_endianswapper_42c2e6ef__1(.endianswapper_42c2e6ef_in(16'h0), 
  .endianswapper_42c2e6ef_out(endianswapper_42c2e6ef_out));
endmodule



module LL1_L_iunzipFilter2D_populateBuffer(CLK, RESET, GO, port_74e37b91_, port_241c8e45_, port_58f1a46c_, port_1a2c8dcf_, RESULT, RESULT_u566, RESULT_u567, RESULT_u568, RESULT_u569, RESULT_u570, RESULT_u571, RESULT_u572, RESULT_u573, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_74e37b91_;
input	[31:0]	port_241c8e45_;
input		port_58f1a46c_;
input	[15:0]	port_1a2c8dcf_;
output		RESULT;
output	[15:0]	RESULT_u566;
output		RESULT_u567;
output	[31:0]	RESULT_u568;
output		RESULT_u569;
output	[31:0]	RESULT_u570;
output	[15:0]	RESULT_u571;
output	[2:0]	RESULT_u572;
output		RESULT_u573;
output		DONE;
wire		simplePinWrite;
wire	[31:0]	add;
wire		and_u1092_u0;
wire		or_u296_u0;
reg		reg_5d954fa8_u0=1'h0;
wire	[31:0]	add_u18;
wire	[15:0]	add_u19;
reg		reg_2e597c75_u0=1'h0;
assign simplePinWrite=GO&{1{GO}};
assign add={port_74e37b91_[15], port_74e37b91_[15], port_74e37b91_[15], port_74e37b91_[15], port_74e37b91_[15], port_74e37b91_[15], port_74e37b91_[15], port_74e37b91_[15], port_74e37b91_[15], port_74e37b91_[15], port_74e37b91_[15], port_74e37b91_[15], port_74e37b91_[15], port_74e37b91_[15], port_74e37b91_[15], port_74e37b91_[15], port_74e37b91_}+32'h0;
assign and_u1092_u0=reg_5d954fa8_u0&port_58f1a46c_;
assign or_u296_u0=and_u1092_u0|RESET;
always @(posedge CLK or posedge GO or posedge or_u296_u0)
begin
if (or_u296_u0)
reg_5d954fa8_u0<=1'h0;
else if (GO)
reg_5d954fa8_u0<=1'h1;
else reg_5d954fa8_u0<=reg_5d954fa8_u0;
end
assign add_u18=port_241c8e45_+32'h1;
assign add_u19=port_74e37b91_+16'h1;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2e597c75_u0<=1'h0;
else reg_2e597c75_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u566=add_u19;
assign RESULT_u567=GO;
assign RESULT_u568=add_u18;
assign RESULT_u569=GO;
assign RESULT_u570=add;
assign RESULT_u571=port_1a2c8dcf_;
assign RESULT_u572=3'h1;
assign RESULT_u573=simplePinWrite;
assign DONE=reg_2e597c75_u0;
endmodule



module LL1_L_iunzipFilter2D_mid1(CLK, RESET, GO, port_60e25201_, port_4fa18e7c_, port_14295d04_, port_1a5e1c20_, port_10388e5c_, port_5ccf9322_, RESULT, RESULT_u574, RESULT_u575, RESULT_u576, RESULT_u577, RESULT_u578, RESULT_u579, RESULT_u580, RESULT_u581, RESULT_u582, RESULT_u583, RESULT_u584, RESULT_u585, RESULT_u586, RESULT_u587, RESULT_u588, RESULT_u589, DONE);
input		CLK;
input		RESET;
input		GO;
input	[31:0]	port_60e25201_;
input	[15:0]	port_4fa18e7c_;
input		port_14295d04_;
input	[15:0]	port_1a5e1c20_;
input		port_10388e5c_;
input	[15:0]	port_5ccf9322_;
output		RESULT;
output	[31:0]	RESULT_u574;
output		RESULT_u575;
output	[15:0]	RESULT_u576;
output		RESULT_u577;
output	[15:0]	RESULT_u578;
output		RESULT_u579;
output	[31:0]	RESULT_u580;
output	[2:0]	RESULT_u581;
output		RESULT_u582;
output	[31:0]	RESULT_u583;
output	[15:0]	RESULT_u584;
output	[2:0]	RESULT_u585;
output	[15:0]	RESULT_u586;
output	[15:0]	RESULT_u587;
output		RESULT_u588;
output		RESULT_u589;
output		DONE;
wire		simplePinWrite;
reg		done_cache_u60=1'h0;
wire		and_u1094_u0;
wire		or_u297_u0;
reg		done_cache_u61_u0=1'h0;
wire		and_u1099_u0;
wire		or_u298_u0;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_538df1a0_instance_RESULT;
wire		and_u1108_u0;
wire		or_u299_u0;
reg		reg_4b6aefd7_u0=1'h0;
wire	[31:0]	add;
wire	[15:0]	add_u20;
wire	[15:0]	simplePinWrite_u173;
wire		simplePinWrite_u174;
wire	[15:0]	simplePinWrite_u175;
reg		reg_0ba433b0_u0=1'h0;
reg		reg_0ba433b0_result_delayed_u0=1'h0;
wire		or_u300_u0;
reg		reg_6d6f405c_u0=1'h0;
reg		reg_0ba433b0_result_delayed_result_delayed_u0=1'h0;
reg	[15:0]	syncEnable_u46=16'h0;
reg		reg_194a1027_u0=1'h0;
reg		reg_6d6f405c_result_delayed_u0=1'h0;
reg	[15:0]	syncEnable_u47_u0=16'h0;
assign simplePinWrite=GO&{1{GO}};
always @(posedge CLK or posedge GO or posedge or_u297_u0)
begin
if (or_u297_u0)
done_cache_u60<=1'h0;
else if (GO)
done_cache_u60<=1'h1;
else done_cache_u60<=done_cache_u60;
end
assign and_u1094_u0=done_cache_u60&port_10388e5c_;
assign or_u297_u0=and_u1094_u0|RESET;
always @(posedge CLK or posedge reg_6d6f405c_result_delayed_u0 or posedge or_u298_u0)
begin
if (or_u298_u0)
done_cache_u61_u0<=1'h0;
else if (reg_6d6f405c_result_delayed_u0)
done_cache_u61_u0<=1'h1;
else done_cache_u61_u0<=done_cache_u61_u0;
end
assign and_u1099_u0=done_cache_u61_u0&port_10388e5c_;
assign or_u298_u0=and_u1099_u0|RESET;
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_538df1a0_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_538df1a0_instance(.GO(reg_194a1027_u0), 
  .port_6062f74a_(syncEnable_u47_u0), .port_77d0cfba_(port_1a5e1c20_), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_538df1a0_instance_RESULT));
assign and_u1108_u0=reg_4b6aefd7_u0&port_10388e5c_;
assign or_u299_u0=and_u1108_u0|RESET;
always @(posedge CLK or posedge reg_0ba433b0_result_delayed_u0 or posedge or_u299_u0)
begin
if (or_u299_u0)
reg_4b6aefd7_u0<=1'h0;
else if (reg_0ba433b0_result_delayed_u0)
reg_4b6aefd7_u0<=1'h1;
else reg_4b6aefd7_u0<=reg_4b6aefd7_u0;
end
assign add=port_60e25201_+32'h1;
assign add_u20=port_4fa18e7c_+16'h1;
assign simplePinWrite_u173=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_538df1a0_instance_RESULT&{16{reg_194a1027_u0}};
assign simplePinWrite_u174=reg_194a1027_u0&{1{reg_194a1027_u0}};
assign simplePinWrite_u175=16'h1&{16{1'h1}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0ba433b0_u0<=1'h0;
else reg_0ba433b0_u0<=reg_194a1027_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0ba433b0_result_delayed_u0<=1'h0;
else reg_0ba433b0_result_delayed_u0<=reg_0ba433b0_u0;
end
assign or_u300_u0=GO|reg_6d6f405c_result_delayed_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6d6f405c_u0<=1'h0;
else reg_6d6f405c_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0ba433b0_result_delayed_result_delayed_u0<=1'h0;
else reg_0ba433b0_result_delayed_result_delayed_u0<=reg_0ba433b0_result_delayed_u0;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u46<=port_5ccf9322_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_194a1027_u0<=1'h0;
else reg_194a1027_u0<=reg_6d6f405c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6d6f405c_result_delayed_u0<=1'h0;
else reg_6d6f405c_result_delayed_u0<=reg_6d6f405c_u0;
end
always @(posedge CLK)
begin
if (reg_6d6f405c_u0)
syncEnable_u47_u0<=port_1a5e1c20_;
end
assign RESULT=GO;
assign RESULT_u574=add;
assign RESULT_u575=GO;
assign RESULT_u576=16'h0;
assign RESULT_u577=GO;
assign RESULT_u578=add_u20;
assign RESULT_u579=or_u300_u0;
assign RESULT_u580=32'h0;
assign RESULT_u581=3'h1;
assign RESULT_u582=reg_0ba433b0_result_delayed_u0;
assign RESULT_u583=32'h0;
assign RESULT_u584=syncEnable_u46;
assign RESULT_u585=3'h1;
assign RESULT_u586=simplePinWrite_u173;
assign RESULT_u587=simplePinWrite_u175;
assign RESULT_u588=simplePinWrite;
assign RESULT_u589=simplePinWrite_u174;
assign DONE=reg_0ba433b0_result_delayed_result_delayed_u0;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_538df1a0_(GO, port_6062f74a_, port_77d0cfba_, RESULT);
input		GO;
input	[15:0]	port_6062f74a_;
input	[15:0]	port_77d0cfba_;
output	[15:0]	RESULT;
wire	[16:0]	add;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_0d6a2ff5_instance_RESULT;
assign add={port_6062f74a_[15], port_6062f74a_}+{port_77d0cfba_[15], port_77d0cfba_};
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_0d6a2ff5_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_0d6a2ff5_instance(.GO(GO), 
  .port_75886818_({add[16], add[16:2]}), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_0d6a2ff5_instance_RESULT));
assign RESULT=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_0d6a2ff5_instance_RESULT;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_0d6a2ff5_(GO, port_75886818_, RESULT);
input		GO;
input	[15:0]	port_75886818_;
output	[15:0]	RESULT;
wire signed	[15:0]	greaterThan_b_signed;
wire		greaterThan;
wire signed	[15:0]	greaterThan_a_signed;
wire		and_u1103_u0;
wire		not_u224_u0;
wire		and_u1104_u0;
wire	[15:0]	mux_u67;
wire		and_u1105_u0;
wire		and_u1106_u0;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_75886818_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign and_u1103_u0=GO&greaterThan;
assign not_u224_u0=~greaterThan;
assign and_u1104_u0=GO&not_u224_u0;
assign mux_u67=(and_u1106_u0)?16'h0:port_75886818_;
assign and_u1105_u0=and_u1104_u0&GO;
assign and_u1106_u0=and_u1103_u0&GO;
assign RESULT=mux_u67;
endmodule



module LL1_L_iunzipFilter2D_midNoConsume1(CLK, RESET, GO, port_60826727_, port_2cb31f5d_, port_09dd1a6b_, RESULT, RESULT_u590, RESULT_u591, RESULT_u592, RESULT_u593, RESULT_u594, RESULT_u595, RESULT_u596, RESULT_u597, RESULT_u598, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_60826727_;
input		port_2cb31f5d_;
input	[15:0]	port_09dd1a6b_;
output		RESULT;
output	[15:0]	RESULT_u590;
output		RESULT_u591;
output	[15:0]	RESULT_u592;
output		RESULT_u593;
output	[31:0]	RESULT_u594;
output	[2:0]	RESULT_u595;
output	[15:0]	RESULT_u596;
output	[15:0]	RESULT_u597;
output		RESULT_u598;
output		DONE;
reg		done_cache_u62=1'h0;
wire		or_u301_u0;
wire		and_u1111_u0;
reg		done_cache_u63_u0=1'h0;
wire		or_u302_u0;
wire		and_u1116_u0;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_799bd57c_instance_RESULT;
wire	[15:0]	add;
wire	[15:0]	simplePinWrite;
wire	[15:0]	simplePinWrite_u176;
wire		simplePinWrite_u177;
reg	[15:0]	syncEnable_u48=16'h0;
wire		or_u303_u0;
reg		reg_5ad40d5f_u0=1'h0;
reg		reg_5ad40d5f_result_delayed_u0=1'h0;
reg		reg_3827c284_u0=1'h0;
reg		reg_5ad40d5f_result_delayed_result_delayed_u0=1'h0;
reg		reg_20368bde_u0=1'h0;
always @(posedge CLK or posedge GO or posedge or_u301_u0)
begin
if (or_u301_u0)
done_cache_u62<=1'h0;
else if (GO)
done_cache_u62<=1'h1;
else done_cache_u62<=done_cache_u62;
end
assign or_u301_u0=and_u1111_u0|RESET;
assign and_u1111_u0=done_cache_u62&port_2cb31f5d_;
always @(posedge CLK or posedge reg_5ad40d5f_u0 or posedge or_u302_u0)
begin
if (or_u302_u0)
done_cache_u63_u0<=1'h0;
else if (reg_5ad40d5f_u0)
done_cache_u63_u0<=1'h1;
else done_cache_u63_u0<=done_cache_u63_u0;
end
assign or_u302_u0=and_u1116_u0|RESET;
assign and_u1116_u0=done_cache_u63_u0&port_2cb31f5d_;
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_799bd57c_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_799bd57c_instance(.GO(reg_5ad40d5f_result_delayed_u0), 
  .port_00f519fd_(port_09dd1a6b_), .port_61373fb2_(syncEnable_u48), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_799bd57c_instance_RESULT));
assign add=port_60826727_+16'h1;
assign simplePinWrite=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_799bd57c_instance_RESULT&{16{reg_5ad40d5f_result_delayed_u0}};
assign simplePinWrite_u176=16'h1&{16{1'h1}};
assign simplePinWrite_u177=reg_5ad40d5f_result_delayed_u0&{1{reg_5ad40d5f_result_delayed_u0}};
always @(posedge CLK)
begin
if (reg_20368bde_u0)
syncEnable_u48<=port_09dd1a6b_;
end
assign or_u303_u0=GO|reg_5ad40d5f_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5ad40d5f_u0<=1'h0;
else reg_5ad40d5f_u0<=reg_20368bde_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5ad40d5f_result_delayed_u0<=1'h0;
else reg_5ad40d5f_result_delayed_u0<=reg_5ad40d5f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3827c284_u0<=1'h0;
else reg_3827c284_u0<=reg_5ad40d5f_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5ad40d5f_result_delayed_result_delayed_u0<=1'h0;
else reg_5ad40d5f_result_delayed_result_delayed_u0<=reg_5ad40d5f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_20368bde_u0<=1'h0;
else reg_20368bde_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u590=16'h0;
assign RESULT_u591=GO;
assign RESULT_u592=add;
assign RESULT_u593=or_u303_u0;
assign RESULT_u594=32'h0;
assign RESULT_u595=3'h1;
assign RESULT_u596=simplePinWrite;
assign RESULT_u597=simplePinWrite_u176;
assign RESULT_u598=simplePinWrite_u177;
assign DONE=reg_3827c284_u0;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_799bd57c_(GO, port_00f519fd_, port_61373fb2_, RESULT);
input		GO;
input	[15:0]	port_00f519fd_;
input	[15:0]	port_61373fb2_;
output	[15:0]	RESULT;
wire	[16:0]	add;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_0a66210c_instance_RESULT;
assign add={port_61373fb2_[15], port_61373fb2_}+{port_00f519fd_[15], port_00f519fd_};
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_0a66210c_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_0a66210c_instance(.GO(GO), 
  .port_012189c0_({add[16], add[16:2]}), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_0a66210c_instance_RESULT));
assign RESULT=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_0a66210c_instance_RESULT;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_0a66210c_(GO, port_012189c0_, RESULT);
input		GO;
input	[15:0]	port_012189c0_;
output	[15:0]	RESULT;
wire signed	[15:0]	greaterThan_a_signed;
wire		greaterThan;
wire signed	[15:0]	greaterThan_b_signed;
wire		and_u1120_u0;
wire		not_u225_u0;
wire		and_u1121_u0;
wire		and_u1122_u0;
wire		and_u1123_u0;
wire	[15:0]	mux_u68;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_012189c0_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign and_u1120_u0=GO&not_u225_u0;
assign not_u225_u0=~greaterThan;
assign and_u1121_u0=GO&greaterThan;
assign and_u1122_u0=and_u1121_u0&GO;
assign and_u1123_u0=and_u1120_u0&GO;
assign mux_u68=(and_u1123_u0)?port_012189c0_:16'h0;
assign RESULT=mux_u68;
endmodule



module LL1_L_iunzipFilter2D_topLeft(CLK, RESET, GO, port_37621793_, port_327d2b21_, port_25f1e81f_, port_2475269b_, port_0b3965ec_, port_4341b031_, port_65941495_, RESULT, RESULT_u599, RESULT_u600, RESULT_u601, RESULT_u602, RESULT_u603, RESULT_u604, RESULT_u605, RESULT_u606, RESULT_u607, RESULT_u608, RESULT_u609, RESULT_u610, RESULT_u611, RESULT_u612, RESULT_u613, RESULT_u614, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_37621793_;
input	[31:0]	port_327d2b21_;
input	[15:0]	port_25f1e81f_;
input		port_2475269b_;
input	[15:0]	port_0b3965ec_;
input		port_4341b031_;
input	[15:0]	port_65941495_;
output		RESULT;
output	[15:0]	RESULT_u599;
output		RESULT_u600;
output	[31:0]	RESULT_u601;
output		RESULT_u602;
output	[15:0]	RESULT_u603;
output		RESULT_u604;
output	[31:0]	RESULT_u605;
output	[2:0]	RESULT_u606;
output		RESULT_u607;
output	[31:0]	RESULT_u608;
output	[15:0]	RESULT_u609;
output	[2:0]	RESULT_u610;
output	[15:0]	RESULT_u611;
output	[15:0]	RESULT_u612;
output		RESULT_u613;
output		RESULT_u614;
output		DONE;
wire		simplePinWrite;
wire		or_u304_u0;
wire		and_u1125_u0;
reg		done_cache_u64=1'h0;
wire		or_u305_u0;
wire		and_u1128_u0;
reg		done_cache_u65_u0=1'h0;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_3b1abe50_instance_RESULT;
wire	[31:0]	add;
reg		reg_5144fbb7_u0=1'h0;
wire		or_u306_u0;
wire		and_u1136_u0;
wire	[15:0]	add_u21;
wire	[31:0]	add_u22;
wire	[15:0]	simplePinWrite_u178;
wire		simplePinWrite_u179;
wire	[15:0]	simplePinWrite_u180;
reg		reg_36881d99_u0=1'h0;
wire	[31:0]	mux_u70;
wire		or_u307_u0;
reg		reg_2c748855_u0=1'h0;
reg		reg_702b0800_u0=1'h0;
reg		reg_2c748855_result_delayed_u0=1'h0;
reg	[15:0]	syncEnable_u49=16'h0;
reg	[31:0]	syncEnable_u50_u0=32'h0;
reg		reg_702b0800_result_delayed_u0=1'h0;
reg	[15:0]	syncEnable_u51_u0=16'h0;
reg		reg_2c748855_result_delayed_result_delayed_u0=1'h0;
assign simplePinWrite=GO&{1{GO}};
assign or_u304_u0=and_u1125_u0|RESET;
assign and_u1125_u0=done_cache_u64&port_4341b031_;
always @(posedge CLK or posedge GO or posedge or_u304_u0)
begin
if (or_u304_u0)
done_cache_u64<=1'h0;
else if (GO)
done_cache_u64<=1'h1;
else done_cache_u64<=done_cache_u64;
end
assign or_u305_u0=and_u1128_u0|RESET;
assign and_u1128_u0=done_cache_u65_u0&port_4341b031_;
always @(posedge CLK or posedge reg_702b0800_result_delayed_u0 or posedge or_u305_u0)
begin
if (or_u305_u0)
done_cache_u65_u0<=1'h0;
else if (reg_702b0800_result_delayed_u0)
done_cache_u65_u0<=1'h1;
else done_cache_u65_u0<=done_cache_u65_u0;
end
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_3b1abe50_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_3b1abe50_instance(.GO(reg_2c748855_u0), 
  .port_241ad0ac_(syncEnable_u51_u0), .port_72dde13c_(port_0b3965ec_), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_3b1abe50_instance_RESULT));
assign add=port_327d2b21_+32'h0;
always @(posedge CLK or posedge reg_2c748855_result_delayed_result_delayed_u0 or posedge or_u306_u0)
begin
if (or_u306_u0)
reg_5144fbb7_u0<=1'h0;
else if (reg_2c748855_result_delayed_result_delayed_u0)
reg_5144fbb7_u0<=1'h1;
else reg_5144fbb7_u0<=reg_5144fbb7_u0;
end
assign or_u306_u0=and_u1136_u0|RESET;
assign and_u1136_u0=reg_5144fbb7_u0&port_4341b031_;
assign add_u21=port_25f1e81f_+16'h1;
assign add_u22=port_327d2b21_+32'h1;
assign simplePinWrite_u178=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_3b1abe50_instance_RESULT&{16{reg_2c748855_u0}};
assign simplePinWrite_u179=reg_2c748855_u0&{1{reg_2c748855_u0}};
assign simplePinWrite_u180=16'h1&{16{1'h1}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_36881d99_u0<=1'h0;
else reg_36881d99_u0<=reg_2c748855_result_delayed_result_delayed_u0;
end
assign mux_u70=({32{reg_2c748855_result_delayed_result_delayed_u0}}&syncEnable_u50_u0)|({32{GO}}&32'h0)|({32{reg_702b0800_result_delayed_u0}}&32'h0);
assign or_u307_u0=GO|reg_702b0800_result_delayed_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2c748855_u0<=1'h0;
else reg_2c748855_u0<=reg_702b0800_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_702b0800_u0<=1'h0;
else reg_702b0800_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2c748855_result_delayed_u0<=1'h0;
else reg_2c748855_result_delayed_u0<=reg_2c748855_u0;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u49<=port_65941495_;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u50_u0<=add;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_702b0800_result_delayed_u0<=1'h0;
else reg_702b0800_result_delayed_u0<=reg_702b0800_u0;
end
always @(posedge CLK)
begin
if (reg_702b0800_u0)
syncEnable_u51_u0<=port_0b3965ec_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2c748855_result_delayed_result_delayed_u0<=1'h0;
else reg_2c748855_result_delayed_result_delayed_u0<=reg_2c748855_result_delayed_u0;
end
assign RESULT=GO;
assign RESULT_u599=16'h0;
assign RESULT_u600=GO;
assign RESULT_u601=add_u22;
assign RESULT_u602=GO;
assign RESULT_u603=add_u21;
assign RESULT_u604=or_u307_u0;
assign RESULT_u605=mux_u70;
assign RESULT_u606=3'h1;
assign RESULT_u607=reg_2c748855_result_delayed_result_delayed_u0;
assign RESULT_u608=mux_u70;
assign RESULT_u609=syncEnable_u49;
assign RESULT_u610=3'h1;
assign RESULT_u611=simplePinWrite_u178;
assign RESULT_u612=simplePinWrite_u180;
assign RESULT_u613=simplePinWrite;
assign RESULT_u614=simplePinWrite_u179;
assign DONE=reg_36881d99_u0;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_3b1abe50_(GO, port_241ad0ac_, port_72dde13c_, RESULT);
input		GO;
input	[15:0]	port_241ad0ac_;
input	[15:0]	port_72dde13c_;
output	[15:0]	RESULT;
wire	[16:0]	add;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_6f963799_instance_RESULT;
assign add={port_241ad0ac_[15], port_241ad0ac_}+{port_72dde13c_[15], port_72dde13c_};
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_6f963799_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_6f963799_instance(.GO(GO), 
  .port_6aa560c4_({add[16], add[16:2]}), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_6f963799_instance_RESULT));
assign RESULT=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_6f963799_instance_RESULT;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_6f963799_(GO, port_6aa560c4_, RESULT);
input		GO;
input	[15:0]	port_6aa560c4_;
output	[15:0]	RESULT;
wire		greaterThan;
wire signed	[15:0]	greaterThan_a_signed;
wire signed	[15:0]	greaterThan_b_signed;
wire		and_u1132_u0;
wire		and_u1133_u0;
wire		not_u226_u0;
wire	[15:0]	mux_u69;
wire		and_u1134_u0;
wire		and_u1135_u0;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_6aa560c4_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign and_u1132_u0=GO&greaterThan;
assign and_u1133_u0=GO&not_u226_u0;
assign not_u226_u0=~greaterThan;
assign mux_u69=(and_u1135_u0)?16'h0:port_6aa560c4_;
assign and_u1134_u0=and_u1133_u0&GO;
assign and_u1135_u0=and_u1132_u0&GO;
assign RESULT=mux_u69;
endmodule



module LL1_L_iunzipFilter2D_donePopulateBuffer(CLK, RESET, GO, RESULT, RESULT_u615, DONE);
input		CLK;
input		RESET;
input		GO;
output		RESULT;
output	[15:0]	RESULT_u615;
output		DONE;
reg		reg_15580b3b_u0=1'h0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_15580b3b_u0<=1'h0;
else reg_15580b3b_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u615=16'h0;
assign DONE=reg_15580b3b_u0;
endmodule



module LL1_L_iunzipFilter2D_bottomRightNoConsume1(CLK, RESET, GO, port_1bf2f003_, port_727877ba_, port_16605d60_, RESULT, RESULT_u616, RESULT_u617, RESULT_u618, RESULT_u619, RESULT_u620, RESULT_u621, RESULT_u622, RESULT_u623, RESULT_u624, RESULT_u625, RESULT_u626, RESULT_u627, RESULT_u628, RESULT_u629, RESULT_u630, DONE);
input		CLK;
input		RESET;
input		GO;
input		port_1bf2f003_;
input		port_727877ba_;
input	[15:0]	port_16605d60_;
output		RESULT;
output	[15:0]	RESULT_u616;
output		RESULT_u617;
output	[15:0]	RESULT_u618;
output		RESULT_u619;
output	[15:0]	RESULT_u620;
output		RESULT_u621;
output	[31:0]	RESULT_u622;
output		RESULT_u623;
output		RESULT_u624;
output		RESULT_u625;
output	[31:0]	RESULT_u626;
output	[2:0]	RESULT_u627;
output	[15:0]	RESULT_u628;
output	[15:0]	RESULT_u629;
output		RESULT_u630;
output		DONE;
wire		and_u1139_u0;
reg		done_cache_u66=1'h0;
wire		or_u308_u0;
wire		and_u1144_u0;
wire		or_u309_u0;
reg		done_cache_u67_u0=1'h0;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_23f12cad_instance_RESULT;
wire		not_u228;
wire	[15:0]	simplePinWrite;
wire		simplePinWrite_u181;
wire	[15:0]	simplePinWrite_u182;
wire		or_u310_u0;
reg		reg_0669d04c_u0=1'h0;
reg	[15:0]	syncEnable_u52=16'h0;
reg		reg_55e061ac_u0=1'h0;
reg		reg_54bfb1f0_u0=1'h0;
reg		reg_0669d04c_result_delayed_u0=1'h0;
reg		reg_54bfb1f0_result_delayed_u0=1'h0;
assign and_u1139_u0=done_cache_u66&port_727877ba_;
always @(posedge CLK or posedge GO or posedge or_u308_u0)
begin
if (or_u308_u0)
done_cache_u66<=1'h0;
else if (GO)
done_cache_u66<=1'h1;
else done_cache_u66<=done_cache_u66;
end
assign or_u308_u0=and_u1139_u0|RESET;
assign and_u1144_u0=done_cache_u67_u0&port_727877ba_;
assign or_u309_u0=and_u1144_u0|RESET;
always @(posedge CLK or posedge reg_54bfb1f0_result_delayed_u0 or posedge or_u309_u0)
begin
if (or_u309_u0)
done_cache_u67_u0<=1'h0;
else if (reg_54bfb1f0_result_delayed_u0)
done_cache_u67_u0<=1'h1;
else done_cache_u67_u0<=done_cache_u67_u0;
end
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_23f12cad_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_23f12cad_instance(.GO(reg_0669d04c_u0), 
  .port_77294153_(syncEnable_u52), .port_2b2800cb_(port_16605d60_), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_23f12cad_instance_RESULT));
assign not_u228=!port_1bf2f003_;
assign simplePinWrite=16'h1&{16{1'h1}};
assign simplePinWrite_u181=reg_0669d04c_u0&{1{reg_0669d04c_u0}};
assign simplePinWrite_u182=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_23f12cad_instance_RESULT&{16{reg_0669d04c_u0}};
assign or_u310_u0=GO|reg_54bfb1f0_result_delayed_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0669d04c_u0<=1'h0;
else reg_0669d04c_u0<=reg_54bfb1f0_result_delayed_u0;
end
always @(posedge CLK)
begin
if (reg_54bfb1f0_u0)
syncEnable_u52<=port_16605d60_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_55e061ac_u0<=1'h0;
else reg_55e061ac_u0<=reg_0669d04c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_54bfb1f0_u0<=1'h0;
else reg_54bfb1f0_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0669d04c_result_delayed_u0<=1'h0;
else reg_0669d04c_result_delayed_u0<=reg_0669d04c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_54bfb1f0_result_delayed_u0<=1'h0;
else reg_54bfb1f0_result_delayed_u0<=reg_54bfb1f0_u0;
end
assign RESULT=GO;
assign RESULT_u616=16'h0;
assign RESULT_u617=GO;
assign RESULT_u618=16'h0;
assign RESULT_u619=GO;
assign RESULT_u620=16'h0;
assign RESULT_u621=GO;
assign RESULT_u622=32'h0;
assign RESULT_u623=GO;
assign RESULT_u624=not_u228;
assign RESULT_u625=or_u310_u0;
assign RESULT_u626=32'h0;
assign RESULT_u627=3'h1;
assign RESULT_u628=simplePinWrite_u182;
assign RESULT_u629=simplePinWrite;
assign RESULT_u630=simplePinWrite_u181;
assign DONE=reg_55e061ac_u0;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_23f12cad_(GO, port_77294153_, port_2b2800cb_, RESULT);
input		GO;
input	[15:0]	port_77294153_;
input	[15:0]	port_2b2800cb_;
output	[15:0]	RESULT;
wire	[16:0]	add;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_5df3fdbb_instance_RESULT;
assign add={port_77294153_[15], port_77294153_}+{port_2b2800cb_[15], port_2b2800cb_};
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_5df3fdbb_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_5df3fdbb_instance(.GO(GO), 
  .port_7bf5c84b_({add[16], add[16:2]}), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_5df3fdbb_instance_RESULT));
assign RESULT=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_5df3fdbb_instance_RESULT;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_5df3fdbb_(GO, port_7bf5c84b_, RESULT);
input		GO;
input	[15:0]	port_7bf5c84b_;
output	[15:0]	RESULT;
wire		greaterThan;
wire signed	[15:0]	greaterThan_b_signed;
wire signed	[15:0]	greaterThan_a_signed;
wire		not_u227_u0;
wire		and_u1148_u0;
wire		and_u1149_u0;
wire		and_u1150_u0;
wire	[15:0]	mux_u71;
wire		and_u1151_u0;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_7bf5c84b_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign not_u227_u0=~greaterThan;
assign and_u1148_u0=GO&greaterThan;
assign and_u1149_u0=GO&not_u227_u0;
assign and_u1150_u0=and_u1149_u0&GO;
assign mux_u71=(and_u1151_u0)?16'h0:port_7bf5c84b_;
assign and_u1151_u0=and_u1148_u0&GO;
assign RESULT=mux_u71;
endmodule



module LL1_L_iunzipFilter2D_mid2(CLK, RESET, GO, port_02e503c9_, port_2ff1ab3b_, port_26472692_, port_160d8dbf_, port_4827c421_, port_564f706b_, RESULT, RESULT_u631, RESULT_u632, RESULT_u633, RESULT_u634, RESULT_u635, RESULT_u636, RESULT_u637, RESULT_u638, RESULT_u639, RESULT_u640, RESULT_u641, RESULT_u642, RESULT_u643, RESULT_u644, RESULT_u645, RESULT_u646, DONE);
input		CLK;
input		RESET;
input		GO;
input	[31:0]	port_02e503c9_;
input	[15:0]	port_2ff1ab3b_;
input		port_26472692_;
input	[15:0]	port_160d8dbf_;
input		port_4827c421_;
input	[15:0]	port_564f706b_;
output		RESULT;
output	[31:0]	RESULT_u631;
output		RESULT_u632;
output	[15:0]	RESULT_u633;
output		RESULT_u634;
output	[15:0]	RESULT_u635;
output		RESULT_u636;
output	[31:0]	RESULT_u637;
output	[2:0]	RESULT_u638;
output		RESULT_u639;
output	[31:0]	RESULT_u640;
output	[15:0]	RESULT_u641;
output	[2:0]	RESULT_u642;
output	[15:0]	RESULT_u643;
output		RESULT_u644;
output	[15:0]	RESULT_u645;
output		RESULT_u646;
output		DONE;
wire		simplePinWrite;
wire		or_u311_u0;
wire		and_u1153_u0;
reg		done_cache_u68=1'h0;
wire		and_u1158_u0;
wire		or_u312_u0;
reg		done_cache_u69_u0=1'h0;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_05e28cb2_instance_RESULT;
wire		or_u313_u0;
reg		reg_34f6fdfd_u0=1'h0;
wire		and_u1167_u0;
wire	[31:0]	add;
wire	[15:0]	add_u23;
wire	[15:0]	simplePinWrite_u183;
wire	[15:0]	simplePinWrite_u184;
wire		simplePinWrite_u185;
reg		reg_7228903b_u0=1'h0;
wire		or_u314_u0;
reg		reg_7228903b_result_delayed_u0=1'h0;
reg		reg_2eaceff9_u0=1'h0;
reg	[15:0]	syncEnable_u53=16'h0;
reg		reg_315986cb_u0=1'h0;
reg		reg_4c8bff13_u0=1'h0;
reg	[15:0]	syncEnable_u54_u0=16'h0;
reg		reg_7228903b_result_delayed_result_delayed_u0=1'h0;
assign simplePinWrite=GO&{1{GO}};
assign or_u311_u0=and_u1153_u0|RESET;
assign and_u1153_u0=done_cache_u68&port_4827c421_;
always @(posedge CLK or posedge GO or posedge or_u311_u0)
begin
if (or_u311_u0)
done_cache_u68<=1'h0;
else if (GO)
done_cache_u68<=1'h1;
else done_cache_u68<=done_cache_u68;
end
assign and_u1158_u0=done_cache_u69_u0&port_4827c421_;
assign or_u312_u0=and_u1158_u0|RESET;
always @(posedge CLK or posedge reg_315986cb_u0 or posedge or_u312_u0)
begin
if (or_u312_u0)
done_cache_u69_u0<=1'h0;
else if (reg_315986cb_u0)
done_cache_u69_u0<=1'h1;
else done_cache_u69_u0<=done_cache_u69_u0;
end
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_05e28cb2_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_05e28cb2_instance(.GO(reg_2eaceff9_u0), 
  .port_52c7e686_(port_160d8dbf_), .port_6c2a9470_(syncEnable_u54_u0), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_05e28cb2_instance_RESULT));
assign or_u313_u0=and_u1167_u0|RESET;
always @(posedge CLK or posedge reg_7228903b_result_delayed_u0 or posedge or_u313_u0)
begin
if (or_u313_u0)
reg_34f6fdfd_u0<=1'h0;
else if (reg_7228903b_result_delayed_u0)
reg_34f6fdfd_u0<=1'h1;
else reg_34f6fdfd_u0<=reg_34f6fdfd_u0;
end
assign and_u1167_u0=reg_34f6fdfd_u0&port_4827c421_;
assign add=port_02e503c9_+32'h1;
assign add_u23=port_2ff1ab3b_+16'h1;
assign simplePinWrite_u183=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_05e28cb2_instance_RESULT&{16{reg_2eaceff9_u0}};
assign simplePinWrite_u184=16'h1&{16{1'h1}};
assign simplePinWrite_u185=reg_2eaceff9_u0&{1{reg_2eaceff9_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7228903b_u0<=1'h0;
else reg_7228903b_u0<=reg_2eaceff9_u0;
end
assign or_u314_u0=GO|reg_315986cb_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7228903b_result_delayed_u0<=1'h0;
else reg_7228903b_result_delayed_u0<=reg_7228903b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2eaceff9_u0<=1'h0;
else reg_2eaceff9_u0<=reg_315986cb_u0;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u53<=port_564f706b_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_315986cb_u0<=1'h0;
else reg_315986cb_u0<=reg_4c8bff13_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4c8bff13_u0<=1'h0;
else reg_4c8bff13_u0<=GO;
end
always @(posedge CLK)
begin
if (reg_4c8bff13_u0)
syncEnable_u54_u0<=port_160d8dbf_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7228903b_result_delayed_result_delayed_u0<=1'h0;
else reg_7228903b_result_delayed_result_delayed_u0<=reg_7228903b_result_delayed_u0;
end
assign RESULT=GO;
assign RESULT_u631=add;
assign RESULT_u632=GO;
assign RESULT_u633=16'h0;
assign RESULT_u634=GO;
assign RESULT_u635=add_u23;
assign RESULT_u636=or_u314_u0;
assign RESULT_u637=32'h0;
assign RESULT_u638=3'h1;
assign RESULT_u639=reg_7228903b_result_delayed_u0;
assign RESULT_u640=32'h0;
assign RESULT_u641=syncEnable_u53;
assign RESULT_u642=3'h1;
assign RESULT_u643=simplePinWrite_u183;
assign RESULT_u644=simplePinWrite;
assign RESULT_u645=simplePinWrite_u184;
assign RESULT_u646=simplePinWrite_u185;
assign DONE=reg_7228903b_result_delayed_result_delayed_u0;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_05e28cb2_(GO, port_52c7e686_, port_6c2a9470_, RESULT);
input		GO;
input	[15:0]	port_52c7e686_;
input	[15:0]	port_6c2a9470_;
output	[15:0]	RESULT;
wire	[15:0]	subtract;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_60bdb814_instance_RESULT;
assign subtract=port_6c2a9470_-port_52c7e686_;
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_60bdb814_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_60bdb814_instance(.GO(GO), 
  .port_7aa2b135_({subtract[15], subtract[15:1]}), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_60bdb814_instance_RESULT));
assign RESULT=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_60bdb814_instance_RESULT;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_60bdb814_(GO, port_7aa2b135_, RESULT);
input		GO;
input	[15:0]	port_7aa2b135_;
output	[15:0]	RESULT;
wire signed	[15:0]	greaterThan_a_signed;
wire signed	[15:0]	greaterThan_b_signed;
wire		greaterThan;
wire		not_u229_u0;
wire		and_u1162_u0;
wire		and_u1163_u0;
wire	[15:0]	mux_u72;
wire		and_u1164_u0;
wire		and_u1165_u0;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_7aa2b135_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign not_u229_u0=~greaterThan;
assign and_u1162_u0=GO&not_u229_u0;
assign and_u1163_u0=GO&greaterThan;
assign mux_u72=(and_u1165_u0)?port_7aa2b135_:16'h0;
assign and_u1164_u0=and_u1163_u0&GO;
assign and_u1165_u0=and_u1162_u0&GO;
assign RESULT=mux_u72;
endmodule



module LL1_L_iunzipFilter2D_midRightNoConsume1(CLK, RESET, GO, port_78715e37_, port_157318c1_, port_7b7c41d3_, port_260281da_, RESULT, RESULT_u647, RESULT_u648, RESULT_u649, RESULT_u650, RESULT_u651, RESULT_u652, RESULT_u653, RESULT_u654, RESULT_u655, RESULT_u656, RESULT_u657, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_78715e37_;
input		port_157318c1_;
input		port_7b7c41d3_;
input	[15:0]	port_260281da_;
output		RESULT;
output	[15:0]	RESULT_u647;
output		RESULT_u648;
output	[15:0]	RESULT_u649;
output		RESULT_u650;
output		RESULT_u651;
output		RESULT_u652;
output	[31:0]	RESULT_u653;
output	[2:0]	RESULT_u654;
output	[15:0]	RESULT_u655;
output	[15:0]	RESULT_u656;
output		RESULT_u657;
output		DONE;
reg		done_cache_u70=1'h0;
wire		and_u1170_u0;
wire		or_u315_u0;
reg		done_cache_u71_u0=1'h0;
wire		and_u1175_u0;
wire		or_u316_u0;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_32b8e3ff_instance_RESULT;
wire	[15:0]	add;
wire		not_u231;
wire	[15:0]	simplePinWrite;
wire	[15:0]	simplePinWrite_u186;
wire		simplePinWrite_u187;
reg	[15:0]	syncEnable_u55=16'h0;
reg		reg_684af871_u0=1'h0;
reg		reg_684af871_result_delayed_u0=1'h0;
reg		reg_01bf3327_u0=1'h0;
reg		reg_18ef5223_u0=1'h0;
wire		or_u317_u0;
reg		reg_01bf3327_result_delayed_u0=1'h0;
always @(posedge CLK or posedge GO or posedge or_u315_u0)
begin
if (or_u315_u0)
done_cache_u70<=1'h0;
else if (GO)
done_cache_u70<=1'h1;
else done_cache_u70<=done_cache_u70;
end
assign and_u1170_u0=done_cache_u70&port_7b7c41d3_;
assign or_u315_u0=and_u1170_u0|RESET;
always @(posedge CLK or posedge reg_01bf3327_result_delayed_u0 or posedge or_u316_u0)
begin
if (or_u316_u0)
done_cache_u71_u0<=1'h0;
else if (reg_01bf3327_result_delayed_u0)
done_cache_u71_u0<=1'h1;
else done_cache_u71_u0<=done_cache_u71_u0;
end
assign and_u1175_u0=done_cache_u71_u0&port_7b7c41d3_;
assign or_u316_u0=and_u1175_u0|RESET;
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_32b8e3ff_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_32b8e3ff_instance(.GO(reg_18ef5223_u0), 
  .port_6b967ae7_(port_260281da_), .port_5394a74f_(syncEnable_u55), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_32b8e3ff_instance_RESULT));
assign add=port_78715e37_+16'h1;
assign not_u231=!port_157318c1_;
assign simplePinWrite=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_32b8e3ff_instance_RESULT&{16{reg_18ef5223_u0}};
assign simplePinWrite_u186=16'h1&{16{1'h1}};
assign simplePinWrite_u187=reg_18ef5223_u0&{1{reg_18ef5223_u0}};
always @(posedge CLK)
begin
if (reg_01bf3327_u0)
syncEnable_u55<=port_260281da_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_684af871_u0<=1'h0;
else reg_684af871_u0<=reg_18ef5223_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_684af871_result_delayed_u0<=1'h0;
else reg_684af871_result_delayed_u0<=reg_684af871_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01bf3327_u0<=1'h0;
else reg_01bf3327_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_18ef5223_u0<=1'h0;
else reg_18ef5223_u0<=reg_01bf3327_result_delayed_u0;
end
assign or_u317_u0=GO|reg_01bf3327_result_delayed_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01bf3327_result_delayed_u0<=1'h0;
else reg_01bf3327_result_delayed_u0<=reg_01bf3327_u0;
end
assign RESULT=GO;
assign RESULT_u647=add;
assign RESULT_u648=GO;
assign RESULT_u649=16'h0;
assign RESULT_u650=GO;
assign RESULT_u651=not_u231;
assign RESULT_u652=or_u317_u0;
assign RESULT_u653=32'h0;
assign RESULT_u654=3'h1;
assign RESULT_u655=simplePinWrite;
assign RESULT_u656=simplePinWrite_u186;
assign RESULT_u657=simplePinWrite_u187;
assign DONE=reg_684af871_result_delayed_u0;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_32b8e3ff_(GO, port_6b967ae7_, port_5394a74f_, RESULT);
input		GO;
input	[15:0]	port_6b967ae7_;
input	[15:0]	port_5394a74f_;
output	[15:0]	RESULT;
wire	[16:0]	add;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_1d1a1cdc_instance_RESULT;
assign add={port_5394a74f_[15], port_5394a74f_}+{port_6b967ae7_[15], port_6b967ae7_};
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_1d1a1cdc_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_1d1a1cdc_instance(.GO(GO), 
  .port_7ccd9fa8_({add[16], add[16:2]}), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_1d1a1cdc_instance_RESULT));
assign RESULT=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_1d1a1cdc_instance_RESULT;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_1d1a1cdc_(GO, port_7ccd9fa8_, RESULT);
input		GO;
input	[15:0]	port_7ccd9fa8_;
output	[15:0]	RESULT;
wire signed	[15:0]	greaterThan_a_signed;
wire signed	[15:0]	greaterThan_b_signed;
wire		greaterThan;
wire		and_u1179_u0;
wire		and_u1180_u0;
wire		not_u230_u0;
wire		and_u1181_u0;
wire	[15:0]	mux_u73;
wire		and_u1182_u0;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_7ccd9fa8_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign and_u1179_u0=GO&not_u230_u0;
assign and_u1180_u0=GO&greaterThan;
assign not_u230_u0=~greaterThan;
assign and_u1181_u0=and_u1180_u0&GO;
assign mux_u73=(and_u1181_u0)?16'h0:port_7ccd9fa8_;
assign and_u1182_u0=and_u1179_u0&GO;
assign RESULT=mux_u73;
endmodule



module LL1_L_iunzipFilter2D_bottomRowNoConsume1(CLK, RESET, GO, port_090c0601_, port_2afc9e1d_, port_0baaff02_, RESULT, RESULT_u658, RESULT_u659, RESULT_u660, RESULT_u661, RESULT_u662, RESULT_u663, RESULT_u664, RESULT_u665, RESULT_u666, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_090c0601_;
input		port_2afc9e1d_;
input	[15:0]	port_0baaff02_;
output		RESULT;
output	[15:0]	RESULT_u658;
output		RESULT_u659;
output	[15:0]	RESULT_u660;
output		RESULT_u661;
output	[31:0]	RESULT_u662;
output	[2:0]	RESULT_u663;
output	[15:0]	RESULT_u664;
output	[15:0]	RESULT_u665;
output		RESULT_u666;
output		DONE;
wire		or_u318_u0;
reg		done_cache_u72=1'h0;
wire		and_u1184_u0;
wire		and_u1189_u0;
reg		done_cache_u73_u0=1'h0;
wire		or_u319_u0;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_6cc82aa4_instance_RESULT;
wire	[15:0]	add;
wire	[15:0]	simplePinWrite;
wire		simplePinWrite_u188;
wire	[15:0]	simplePinWrite_u189;
reg		reg_62ed9e80_u0=1'h0;
wire		or_u320_u0;
reg	[15:0]	syncEnable_u56=16'h0;
reg		reg_1eca9562_u0=1'h0;
reg		reg_1eca9562_result_delayed_u0=1'h0;
reg		reg_0ff2022a_u0=1'h0;
reg		reg_62ed9e80_result_delayed_u0=1'h0;
assign or_u318_u0=and_u1184_u0|RESET;
always @(posedge CLK or posedge GO or posedge or_u318_u0)
begin
if (or_u318_u0)
done_cache_u72<=1'h0;
else if (GO)
done_cache_u72<=1'h1;
else done_cache_u72<=done_cache_u72;
end
assign and_u1184_u0=done_cache_u72&port_2afc9e1d_;
assign and_u1189_u0=done_cache_u73_u0&port_2afc9e1d_;
always @(posedge CLK or posedge reg_62ed9e80_result_delayed_u0 or posedge or_u319_u0)
begin
if (or_u319_u0)
done_cache_u73_u0<=1'h0;
else if (reg_62ed9e80_result_delayed_u0)
done_cache_u73_u0<=1'h1;
else done_cache_u73_u0<=done_cache_u73_u0;
end
assign or_u319_u0=and_u1189_u0|RESET;
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_6cc82aa4_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_6cc82aa4_instance(.GO(reg_0ff2022a_u0), 
  .port_0e0fac7a_(syncEnable_u56), .port_3ea0767e_(port_0baaff02_), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_6cc82aa4_instance_RESULT));
assign add=port_090c0601_+16'h1;
assign simplePinWrite=16'h1&{16{1'h1}};
assign simplePinWrite_u188=reg_0ff2022a_u0&{1{reg_0ff2022a_u0}};
assign simplePinWrite_u189=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_6cc82aa4_instance_RESULT&{16{reg_0ff2022a_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_62ed9e80_u0<=1'h0;
else reg_62ed9e80_u0<=GO;
end
assign or_u320_u0=GO|reg_62ed9e80_result_delayed_u0;
always @(posedge CLK)
begin
if (reg_62ed9e80_u0)
syncEnable_u56<=port_0baaff02_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1eca9562_u0<=1'h0;
else reg_1eca9562_u0<=reg_0ff2022a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1eca9562_result_delayed_u0<=1'h0;
else reg_1eca9562_result_delayed_u0<=reg_1eca9562_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0ff2022a_u0<=1'h0;
else reg_0ff2022a_u0<=reg_62ed9e80_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_62ed9e80_result_delayed_u0<=1'h0;
else reg_62ed9e80_result_delayed_u0<=reg_62ed9e80_u0;
end
assign RESULT=GO;
assign RESULT_u658=16'h0;
assign RESULT_u659=GO;
assign RESULT_u660=add;
assign RESULT_u661=or_u320_u0;
assign RESULT_u662=32'h0;
assign RESULT_u663=3'h1;
assign RESULT_u664=simplePinWrite_u189;
assign RESULT_u665=simplePinWrite;
assign RESULT_u666=simplePinWrite_u188;
assign DONE=reg_1eca9562_result_delayed_u0;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_6cc82aa4_(GO, port_0e0fac7a_, port_3ea0767e_, RESULT);
input		GO;
input	[15:0]	port_0e0fac7a_;
input	[15:0]	port_3ea0767e_;
output	[15:0]	RESULT;
wire	[16:0]	add;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_0109403f_instance_RESULT;
assign add={port_0e0fac7a_[15], port_0e0fac7a_}+{port_3ea0767e_[15], port_3ea0767e_};
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_0109403f_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_0109403f_instance(.GO(GO), 
  .port_3454eeda_({add[16], add[16:2]}), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_0109403f_instance_RESULT));
assign RESULT=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_0109403f_instance_RESULT;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_0109403f_(GO, port_3454eeda_, RESULT);
input		GO;
input	[15:0]	port_3454eeda_;
output	[15:0]	RESULT;
wire signed	[15:0]	greaterThan_b_signed;
wire signed	[15:0]	greaterThan_a_signed;
wire		greaterThan;
wire		and_u1193_u0;
wire		not_u232_u0;
wire		and_u1194_u0;
wire		and_u1195_u0;
wire	[15:0]	mux_u74;
wire		and_u1196_u0;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_3454eeda_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign and_u1193_u0=GO&not_u232_u0;
assign not_u232_u0=~greaterThan;
assign and_u1194_u0=GO&greaterThan;
assign and_u1195_u0=and_u1194_u0&GO;
assign mux_u74=(and_u1195_u0)?16'h0:port_3454eeda_;
assign and_u1196_u0=and_u1193_u0&GO;
assign RESULT=mux_u74;
endmodule



module LL1_L_iunzipFilter2D_Kicker_15(CLK, RESET, bus_1e59a7e8_);
input		CLK;
input		RESET;
output		bus_1e59a7e8_;
reg		kicker_2=1'h0;
wire		bus_1a6a6284_;
wire		bus_484f7ad0_;
wire		bus_32d83335_;
reg		kicker_1=1'h0;
wire		bus_65db3e8c_;
reg		kicker_res=1'h0;
always @(posedge CLK)
begin
kicker_2<=bus_32d83335_;
end
assign bus_1a6a6284_=kicker_1&bus_484f7ad0_&bus_65db3e8c_;
assign bus_484f7ad0_=~RESET;
assign bus_32d83335_=bus_484f7ad0_&kicker_1;
always @(posedge CLK)
begin
kicker_1<=bus_484f7ad0_;
end
assign bus_65db3e8c_=~kicker_2;
always @(posedge CLK)
begin
kicker_res<=bus_1a6a6284_;
end
assign bus_1e59a7e8_=kicker_res;
endmodule



module LL1_L_iunzipFilter2D_simplememoryreferee_570ba99f_(bus_24dbf5d8_, bus_1e68ee92_, bus_42b63aee_, bus_4d929d8d_, bus_0dc704d1_, bus_35b4734c_, bus_3ff68fd8_, bus_2e8e26fe_, bus_123b1c5f_, bus_4b4b39e6_, bus_58ff9411_, bus_62c5dd82_, bus_31fab083_, bus_33af7415_);
input		bus_24dbf5d8_;
input		bus_1e68ee92_;
input		bus_42b63aee_;
input	[15:0]	bus_4d929d8d_;
input		bus_0dc704d1_;
input	[15:0]	bus_35b4734c_;
input	[31:0]	bus_3ff68fd8_;
input	[2:0]	bus_2e8e26fe_;
output	[15:0]	bus_123b1c5f_;
output	[31:0]	bus_4b4b39e6_;
output		bus_58ff9411_;
output		bus_62c5dd82_;
output	[2:0]	bus_31fab083_;
output		bus_33af7415_;
assign bus_123b1c5f_=bus_35b4734c_;
assign bus_4b4b39e6_=bus_3ff68fd8_;
assign bus_58ff9411_=bus_0dc704d1_;
assign bus_62c5dd82_=bus_0dc704d1_;
assign bus_31fab083_=3'h1;
assign bus_33af7415_=bus_42b63aee_;
endmodule



module LL1_L_iunzipFilter2D_bottomRowNoConsume2(CLK, RESET, GO, port_72d40a34_, port_2dfef218_, port_1cd6730f_, RESULT, RESULT_u667, RESULT_u668, RESULT_u669, RESULT_u670, RESULT_u671, RESULT_u672, RESULT_u673, RESULT_u674, RESULT_u675, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_72d40a34_;
input		port_2dfef218_;
input	[15:0]	port_1cd6730f_;
output		RESULT;
output	[15:0]	RESULT_u667;
output		RESULT_u668;
output	[15:0]	RESULT_u669;
output		RESULT_u670;
output	[31:0]	RESULT_u671;
output	[2:0]	RESULT_u672;
output	[15:0]	RESULT_u673;
output		RESULT_u674;
output	[15:0]	RESULT_u675;
output		DONE;
reg		done_cache_u74=1'h0;
wire		and_u1199_u0;
wire		or_u321_u0;
wire		or_u322_u0;
wire		and_u1204_u0;
reg		done_cache_u75_u0=1'h0;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_77568265_instance_RESULT;
wire	[15:0]	add;
wire		simplePinWrite;
wire	[15:0]	simplePinWrite_u190;
wire	[15:0]	simplePinWrite_u191;
reg		reg_24ed56f6_u0=1'h0;
wire		or_u323_u0;
reg		reg_5033f266_u0=1'h0;
reg	[15:0]	syncEnable_u57=16'h0;
reg		reg_3a1883a9_u0=1'h0;
reg		reg_6be62207_u0=1'h0;
reg		reg_24ed56f6_result_delayed_u0=1'h0;
always @(posedge CLK or posedge GO or posedge or_u321_u0)
begin
if (or_u321_u0)
done_cache_u74<=1'h0;
else if (GO)
done_cache_u74<=1'h1;
else done_cache_u74<=done_cache_u74;
end
assign and_u1199_u0=done_cache_u74&port_2dfef218_;
assign or_u321_u0=and_u1199_u0|RESET;
assign or_u322_u0=and_u1204_u0|RESET;
assign and_u1204_u0=done_cache_u75_u0&port_2dfef218_;
always @(posedge CLK or posedge reg_3a1883a9_u0 or posedge or_u322_u0)
begin
if (or_u322_u0)
done_cache_u75_u0<=1'h0;
else if (reg_3a1883a9_u0)
done_cache_u75_u0<=1'h1;
else done_cache_u75_u0<=done_cache_u75_u0;
end
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_77568265_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_77568265_instance(.GO(reg_5033f266_u0), 
  .port_375e3c95_(syncEnable_u57), .port_187faf8b_(port_1cd6730f_), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_77568265_instance_RESULT));
assign add=port_72d40a34_+16'h1;
assign simplePinWrite=reg_5033f266_u0&{1{reg_5033f266_u0}};
assign simplePinWrite_u190=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_77568265_instance_RESULT&{16{reg_5033f266_u0}};
assign simplePinWrite_u191=16'h1&{16{1'h1}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_24ed56f6_u0<=1'h0;
else reg_24ed56f6_u0<=reg_5033f266_u0;
end
assign or_u323_u0=GO|reg_3a1883a9_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5033f266_u0<=1'h0;
else reg_5033f266_u0<=reg_3a1883a9_u0;
end
always @(posedge CLK)
begin
if (reg_6be62207_u0)
syncEnable_u57<=port_1cd6730f_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3a1883a9_u0<=1'h0;
else reg_3a1883a9_u0<=reg_6be62207_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6be62207_u0<=1'h0;
else reg_6be62207_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_24ed56f6_result_delayed_u0<=1'h0;
else reg_24ed56f6_result_delayed_u0<=reg_24ed56f6_u0;
end
assign RESULT=GO;
assign RESULT_u667=16'h0;
assign RESULT_u668=GO;
assign RESULT_u669=add;
assign RESULT_u670=or_u323_u0;
assign RESULT_u671=32'h0;
assign RESULT_u672=3'h1;
assign RESULT_u673=simplePinWrite_u190;
assign RESULT_u674=simplePinWrite;
assign RESULT_u675=simplePinWrite_u191;
assign DONE=reg_24ed56f6_result_delayed_u0;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_77568265_(GO, port_375e3c95_, port_187faf8b_, RESULT);
input		GO;
input	[15:0]	port_375e3c95_;
input	[15:0]	port_187faf8b_;
output	[15:0]	RESULT;
wire	[15:0]	subtract;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_0619f7d2_instance_RESULT;
assign subtract=port_375e3c95_-port_187faf8b_;
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_0619f7d2_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_0619f7d2_instance(.GO(GO), 
  .port_46890aea_({subtract[15], subtract[15:1]}), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_0619f7d2_instance_RESULT));
assign RESULT=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_0619f7d2_instance_RESULT;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_0619f7d2_(GO, port_46890aea_, RESULT);
input		GO;
input	[15:0]	port_46890aea_;
output	[15:0]	RESULT;
wire		greaterThan;
wire signed	[15:0]	greaterThan_a_signed;
wire signed	[15:0]	greaterThan_b_signed;
wire		and_u1208_u0;
wire		and_u1209_u0;
wire		not_u233_u0;
wire		and_u1210_u0;
wire	[15:0]	mux_u75;
wire		and_u1211_u0;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_46890aea_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign and_u1208_u0=GO&greaterThan;
assign and_u1209_u0=GO&not_u233_u0;
assign not_u233_u0=~greaterThan;
assign and_u1210_u0=and_u1208_u0&GO;
assign mux_u75=(and_u1210_u0)?16'h0:port_46890aea_;
assign and_u1211_u0=and_u1209_u0&GO;
assign RESULT=mux_u75;
endmodule



module LL1_L_iunzipFilter2D_forge_memory_515x16_3(CLK, ENA, WEA, DINA, ENB, WEB, DINB, ADDRA, ADDRB, DOUTA, DOUTB, DONEA, DONEB);
input		CLK;
input		ENA;
input		WEA;
input	[15:0]	DINA;
input		ENB;
input		WEB;
input	[15:0]	DINB;
input	[31:0]	ADDRA;
input	[31:0]	ADDRB;
output	[15:0]	DOUTA;
output	[15:0]	DOUTB;
output		DONEA;
output		DONEB;
wire		wea_0;
wire		web_0;
wire	[15:0]	pre_douta_0;
wire	[15:0]	pre_doutb_0;
wire	[1:0]	extrasa_0;
wire	[1:0]	extrasb_0;
reg	[15:0]	mux_outa;
reg	[15:0]	mux_outb;
reg	[31:0]	ADDRA_reg;
reg	[31:0]	ADDRB_reg;
reg		rea_done;
reg		wea_done;
reg		web_done;
reg		reb_done;
assign wea_0=WEA&(ADDRA[31:10]==22'h0);
assign web_0=WEB&(ADDRB[31:10]==22'h0);
always @(posedge CLK)
begin
ADDRA_reg<=ADDRA;
end
always @(pre_douta_0)
begin
mux_outa<=pre_douta_0;
end
always @(posedge CLK)
begin
ADDRB_reg<=ADDRB;
end
always @(pre_doutb_0)
begin
mux_outb<=pre_doutb_0;
end
always @(posedge CLK)
begin
wea_done<=WEA;
rea_done<=ENA;
web_done<=WEB;
reb_done<=ENB;
end
assign DONEA=wea_done|rea_done;
assign DONEB=web_done|reb_done;
assign DOUTA=mux_outa;
assign DOUTB=mux_outb;
// Memory array element: COL: 0, ROW: 0
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S18_S18#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S18_S18_instance_1(.CLKA(CLK), 
  .WEA(wea_0), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[15:0]), .DOA(pre_douta_0[15:0]), 
  .DIPA(2'b0), .DOPA(), .CLKB(CLK), .WEB(web_0), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), 
  .DIB(DINB[15:0]), .DOB(pre_doutb_0[15:0]), .DIPB(2'b0), .DOPB());
endmodule



module LL1_L_iunzipFilter2D_structuralmemory_01e37556_(CLK_u1, bus_5916951f_, bus_7f082c33_, bus_2219040d_, bus_4d72aca4_, bus_6b921393_, bus_1b1b36f0_, bus_75697e3b_, bus_369fe81a_, bus_0986c750_, bus_339c133a_, bus_4db85e66_, bus_0189de6b_, bus_44ef805d_, bus_75e069b0_, bus_3e990c66_);
input		CLK_u1;
input		bus_5916951f_;
input	[31:0]	bus_7f082c33_;
input	[2:0]	bus_2219040d_;
input		bus_4d72aca4_;
input		bus_6b921393_;
input	[15:0]	bus_1b1b36f0_;
input	[31:0]	bus_75697e3b_;
input	[2:0]	bus_369fe81a_;
input		bus_0986c750_;
input		bus_339c133a_;
input	[15:0]	bus_4db85e66_;
output	[15:0]	bus_0189de6b_;
output		bus_44ef805d_;
output	[15:0]	bus_75e069b0_;
output		bus_3e990c66_;
wire	[15:0]	bus_7442309c_;
wire	[15:0]	bus_26f6e502_;
wire		or_273dba2e_u0;
reg		logicalMem_69d35e5d_re_delay0_u0=1'h0;
reg		logicalMem_69d35e5d_we_delay0_u0=1'h0;
wire		or_0ab27652_u0;
reg		logicalMem_69d35e5d_re_delay0_u1_u0=1'h0;
wire		or_63c64eb4_u0;
wire		or_1a1769e3_u0;
reg		logicalMem_69d35e5d_we_delay0_u1_u0=1'h0;
LL1_L_iunzipFilter2D_forge_memory_515x16_3 LL1_L_iunzipFilter2D_forge_memory_515x16_3_instance0(.CLK(CLK_u1), 
  .ENA(or_0ab27652_u0), .WEA(bus_6b921393_), .DINA(bus_1b1b36f0_), .ADDRA(bus_7f082c33_), 
  .DOUTA(bus_26f6e502_), .DONEA(), .ENB(or_273dba2e_u0), .WEB(bus_339c133a_), .DINB(bus_4db85e66_), 
  .ADDRB(bus_75697e3b_), .DOUTB(bus_7442309c_), .DONEB());
assign or_273dba2e_u0=bus_0986c750_|bus_339c133a_;
always @(posedge CLK_u1 or posedge bus_5916951f_)
begin
if (bus_5916951f_)
logicalMem_69d35e5d_re_delay0_u0<=1'h0;
else logicalMem_69d35e5d_re_delay0_u0<=bus_0986c750_;
end
always @(posedge CLK_u1 or posedge bus_5916951f_)
begin
if (bus_5916951f_)
logicalMem_69d35e5d_we_delay0_u0<=1'h0;
else logicalMem_69d35e5d_we_delay0_u0<=bus_6b921393_;
end
assign or_0ab27652_u0=bus_4d72aca4_|bus_6b921393_;
always @(posedge CLK_u1 or posedge bus_5916951f_)
begin
if (bus_5916951f_)
logicalMem_69d35e5d_re_delay0_u1_u0<=1'h0;
else logicalMem_69d35e5d_re_delay0_u1_u0<=bus_4d72aca4_;
end
assign or_63c64eb4_u0=logicalMem_69d35e5d_re_delay0_u0|logicalMem_69d35e5d_we_delay0_u1_u0;
assign or_1a1769e3_u0=logicalMem_69d35e5d_re_delay0_u1_u0|logicalMem_69d35e5d_we_delay0_u0;
assign bus_0189de6b_=bus_26f6e502_;
assign bus_44ef805d_=or_1a1769e3_u0;
assign bus_75e069b0_=bus_7442309c_;
assign bus_3e990c66_=or_63c64eb4_u0;
always @(posedge CLK_u1 or posedge bus_5916951f_)
begin
if (bus_5916951f_)
logicalMem_69d35e5d_we_delay0_u1_u0<=1'h0;
else logicalMem_69d35e5d_we_delay0_u1_u0<=bus_339c133a_;
end
endmodule



module LL1_L_iunzipFilter2D_bottomRightNoConsume2(CLK, RESET, GO, port_6ecd2cdc_, port_0eaeaa28_, port_3ee0a27c_, RESULT, RESULT_u676, RESULT_u677, RESULT_u678, RESULT_u679, RESULT_u680, RESULT_u681, RESULT_u682, RESULT_u683, RESULT_u684, RESULT_u685, RESULT_u686, RESULT_u687, RESULT_u688, RESULT_u689, RESULT_u690, DONE);
input		CLK;
input		RESET;
input		GO;
input		port_6ecd2cdc_;
input		port_0eaeaa28_;
input	[15:0]	port_3ee0a27c_;
output		RESULT;
output	[15:0]	RESULT_u676;
output		RESULT_u677;
output	[15:0]	RESULT_u678;
output		RESULT_u679;
output	[15:0]	RESULT_u680;
output		RESULT_u681;
output	[31:0]	RESULT_u682;
output		RESULT_u683;
output		RESULT_u684;
output		RESULT_u685;
output	[31:0]	RESULT_u686;
output	[2:0]	RESULT_u687;
output	[15:0]	RESULT_u688;
output		RESULT_u689;
output	[15:0]	RESULT_u690;
output		DONE;
reg		done_cache_u76=1'h0;
wire		or_u324_u0;
wire		and_u1214_u0;
wire		and_u1219_u0;
wire		or_u325_u0;
reg		done_cache_u77_u0=1'h0;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_59ec89db_instance_RESULT;
wire		not_u235;
wire		simplePinWrite;
wire	[15:0]	simplePinWrite_u192;
wire	[15:0]	simplePinWrite_u193;
reg		reg_4a057739_u0=1'h0;
reg		reg_15b4e4f6_u0=1'h0;
reg		reg_4a057739_result_delayed_u0=1'h0;
reg		reg_155bc105_u0=1'h0;
reg		reg_79c6b34c_u0=1'h0;
reg	[15:0]	syncEnable_u58=16'h0;
wire		or_u326_u0;
always @(posedge CLK or posedge GO or posedge or_u324_u0)
begin
if (or_u324_u0)
done_cache_u76<=1'h0;
else if (GO)
done_cache_u76<=1'h1;
else done_cache_u76<=done_cache_u76;
end
assign or_u324_u0=and_u1214_u0|RESET;
assign and_u1214_u0=done_cache_u76&port_0eaeaa28_;
assign and_u1219_u0=done_cache_u77_u0&port_0eaeaa28_;
assign or_u325_u0=and_u1219_u0|RESET;
always @(posedge CLK or posedge reg_155bc105_u0 or posedge or_u325_u0)
begin
if (or_u325_u0)
done_cache_u77_u0<=1'h0;
else if (reg_155bc105_u0)
done_cache_u77_u0<=1'h1;
else done_cache_u77_u0<=done_cache_u77_u0;
end
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_59ec89db_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_59ec89db_instance(.GO(reg_4a057739_u0), 
  .port_0b5b273c_(syncEnable_u58), .port_3e17bcdb_(port_3ee0a27c_), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_59ec89db_instance_RESULT));
assign not_u235=!port_6ecd2cdc_;
assign simplePinWrite=reg_4a057739_u0&{1{reg_4a057739_u0}};
assign simplePinWrite_u192=16'h1&{16{1'h1}};
assign simplePinWrite_u193=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_59ec89db_instance_RESULT&{16{reg_4a057739_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4a057739_u0<=1'h0;
else reg_4a057739_u0<=reg_155bc105_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_15b4e4f6_u0<=1'h0;
else reg_15b4e4f6_u0<=reg_4a057739_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4a057739_result_delayed_u0<=1'h0;
else reg_4a057739_result_delayed_u0<=reg_4a057739_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_155bc105_u0<=1'h0;
else reg_155bc105_u0<=reg_79c6b34c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_79c6b34c_u0<=1'h0;
else reg_79c6b34c_u0<=GO;
end
always @(posedge CLK)
begin
if (reg_79c6b34c_u0)
syncEnable_u58<=port_3ee0a27c_;
end
assign or_u326_u0=GO|reg_155bc105_u0;
assign RESULT=GO;
assign RESULT_u676=16'h0;
assign RESULT_u677=GO;
assign RESULT_u678=16'h0;
assign RESULT_u679=GO;
assign RESULT_u680=16'h0;
assign RESULT_u681=GO;
assign RESULT_u682=32'h0;
assign RESULT_u683=GO;
assign RESULT_u684=not_u235;
assign RESULT_u685=or_u326_u0;
assign RESULT_u686=32'h0;
assign RESULT_u687=3'h1;
assign RESULT_u688=simplePinWrite_u193;
assign RESULT_u689=simplePinWrite;
assign RESULT_u690=simplePinWrite_u192;
assign DONE=reg_15b4e4f6_u0;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_59ec89db_(GO, port_0b5b273c_, port_3e17bcdb_, RESULT);
input		GO;
input	[15:0]	port_0b5b273c_;
input	[15:0]	port_3e17bcdb_;
output	[15:0]	RESULT;
wire	[15:0]	subtract;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_45395689_instance_RESULT;
assign subtract=port_0b5b273c_-port_3e17bcdb_;
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_45395689_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_45395689_instance(.GO(GO), 
  .port_66a271c4_({subtract[15], subtract[15:1]}), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_45395689_instance_RESULT));
assign RESULT=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_45395689_instance_RESULT;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_45395689_(GO, port_66a271c4_, RESULT);
input		GO;
input	[15:0]	port_66a271c4_;
output	[15:0]	RESULT;
wire signed	[15:0]	greaterThan_a_signed;
wire		greaterThan;
wire signed	[15:0]	greaterThan_b_signed;
wire		and_u1223_u0;
wire		not_u234_u0;
wire		and_u1224_u0;
wire		and_u1225_u0;
wire		and_u1226_u0;
wire	[15:0]	mux_u76;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_66a271c4_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign and_u1223_u0=GO&greaterThan;
assign not_u234_u0=~greaterThan;
assign and_u1224_u0=GO&not_u234_u0;
assign and_u1225_u0=and_u1224_u0&GO;
assign and_u1226_u0=and_u1223_u0&GO;
assign mux_u76=(and_u1226_u0)?16'h0:port_66a271c4_;
assign RESULT=mux_u76;
endmodule



module LL1_L_iunzipFilter2D_endianswapper_38835f81_(endianswapper_38835f81_in, endianswapper_38835f81_out);
input	[15:0]	endianswapper_38835f81_in;
output	[15:0]	endianswapper_38835f81_out;
assign endianswapper_38835f81_out=endianswapper_38835f81_in;
endmodule



module LL1_L_iunzipFilter2D_endianswapper_17bc34ff_(endianswapper_17bc34ff_in, endianswapper_17bc34ff_out);
input	[15:0]	endianswapper_17bc34ff_in;
output	[15:0]	endianswapper_17bc34ff_out;
assign endianswapper_17bc34ff_out=endianswapper_17bc34ff_in;
endmodule



module LL1_L_iunzipFilter2D_stateVar_midPtr(bus_38bd42c5_, bus_00f33b37_, bus_53c01961_, bus_188a6b35_, bus_16d1222c_, bus_122af5f2_, bus_01f7a039_, bus_0aba6433_, bus_698b642e_, bus_2bc2559e_, bus_43c76f68_, bus_0903fe04_, bus_7e6c4fd8_, bus_7955a617_, bus_2551f507_, bus_1a0acc16_, bus_723ff3dc_, bus_2d47447b_, bus_1ed9e97d_, bus_62513a6e_, bus_0a10bc57_, bus_02599f9e_, bus_4f97ace6_, bus_6a732550_, bus_0a1ca6cd_, bus_1a147c05_, bus_7becdf00_, bus_5fec891a_, bus_1fdda57d_, bus_4b200500_, bus_1826a746_, bus_5ce7e0b1_, bus_0b07ce99_, bus_58e8f3e2_, bus_79009f57_, bus_1603d043_, bus_10233de4_, bus_4bb9035f_, bus_087b7bab_, bus_4abfcc53_, bus_6d53b8af_, bus_6c7eeb69_, bus_13e6efa8_, bus_6b6720f0_, bus_7da5ce18_);
input		bus_38bd42c5_;
input		bus_00f33b37_;
input		bus_53c01961_;
input	[15:0]	bus_188a6b35_;
input		bus_16d1222c_;
input	[15:0]	bus_122af5f2_;
input		bus_01f7a039_;
input	[15:0]	bus_0aba6433_;
input		bus_698b642e_;
input	[15:0]	bus_2bc2559e_;
input		bus_43c76f68_;
input	[15:0]	bus_0903fe04_;
input		bus_7e6c4fd8_;
input	[15:0]	bus_7955a617_;
input		bus_2551f507_;
input	[15:0]	bus_1a0acc16_;
input		bus_723ff3dc_;
input	[15:0]	bus_2d47447b_;
input		bus_1ed9e97d_;
input	[15:0]	bus_62513a6e_;
input		bus_0a10bc57_;
input	[15:0]	bus_02599f9e_;
input		bus_4f97ace6_;
input	[15:0]	bus_6a732550_;
input		bus_0a1ca6cd_;
input	[15:0]	bus_1a147c05_;
input		bus_7becdf00_;
input	[15:0]	bus_5fec891a_;
input		bus_1fdda57d_;
input	[15:0]	bus_4b200500_;
input		bus_1826a746_;
input	[15:0]	bus_5ce7e0b1_;
input		bus_0b07ce99_;
input	[15:0]	bus_58e8f3e2_;
input		bus_79009f57_;
input	[15:0]	bus_1603d043_;
input		bus_10233de4_;
input	[15:0]	bus_4bb9035f_;
input		bus_087b7bab_;
input	[15:0]	bus_4abfcc53_;
input		bus_6d53b8af_;
input	[15:0]	bus_6c7eeb69_;
input		bus_13e6efa8_;
input	[15:0]	bus_6b6720f0_;
output	[15:0]	bus_7da5ce18_;
wire	[15:0]	endianswapper_38835f81_out;
wire	[15:0]	endianswapper_17bc34ff_out;
wire		or_37a8df11_u0;
reg	[15:0]	stateVar_midPtr_u1=16'h0;
wire	[15:0]	mux_2dd201ce_u0;
LL1_L_iunzipFilter2D_endianswapper_38835f81_ LL1_L_iunzipFilter2D_endianswapper_38835f81__1(.endianswapper_38835f81_in(stateVar_midPtr_u1), 
  .endianswapper_38835f81_out(endianswapper_38835f81_out));
LL1_L_iunzipFilter2D_endianswapper_17bc34ff_ LL1_L_iunzipFilter2D_endianswapper_17bc34ff__1(.endianswapper_17bc34ff_in(mux_2dd201ce_u0), 
  .endianswapper_17bc34ff_out(endianswapper_17bc34ff_out));
assign bus_7da5ce18_=endianswapper_38835f81_out;
assign or_37a8df11_u0=bus_53c01961_|bus_16d1222c_|bus_01f7a039_|bus_698b642e_|bus_43c76f68_|bus_7e6c4fd8_|bus_2551f507_|bus_723ff3dc_|bus_1ed9e97d_|bus_0a10bc57_|bus_4f97ace6_|bus_0a1ca6cd_|bus_7becdf00_|bus_1fdda57d_|bus_1826a746_|bus_0b07ce99_|bus_79009f57_|bus_10233de4_|bus_087b7bab_|bus_6d53b8af_|bus_13e6efa8_;
always @(posedge bus_38bd42c5_ or posedge bus_00f33b37_)
begin
if (bus_00f33b37_)
stateVar_midPtr_u1<=16'h0;
else if (or_37a8df11_u0)
stateVar_midPtr_u1<=endianswapper_17bc34ff_out;
end
assign mux_2dd201ce_u0=({16{bus_53c01961_}}&bus_188a6b35_)|({16{bus_16d1222c_}}&bus_122af5f2_)|({16{bus_01f7a039_}}&16'h0)|({16{bus_698b642e_}}&bus_2bc2559e_)|({16{bus_43c76f68_}}&bus_0903fe04_)|({16{bus_7e6c4fd8_}}&bus_7955a617_)|({16{bus_2551f507_}}&bus_1a0acc16_)|({16{bus_723ff3dc_}}&bus_2d47447b_)|({16{bus_1ed9e97d_}}&bus_62513a6e_)|({16{bus_0a10bc57_}}&bus_02599f9e_)|({16{bus_4f97ace6_}}&bus_6a732550_)|({16{bus_0a1ca6cd_}}&16'h0)|({16{bus_7becdf00_}}&16'h0)|({16{bus_1fdda57d_}}&16'h0)|({16{bus_1826a746_}}&16'h0)|({16{bus_0b07ce99_}}&bus_58e8f3e2_)|({16{bus_79009f57_}}&bus_1603d043_)|({16{bus_10233de4_}}&bus_4bb9035f_)|({16{bus_087b7bab_}}&bus_4abfcc53_)|({16{bus_6d53b8af_}}&16'h0)|({16{bus_13e6efa8_}}&16'h0);
endmodule



module LL1_L_iunzipFilter2D_endianswapper_717afd68_(endianswapper_717afd68_in, endianswapper_717afd68_out);
input	[15:0]	endianswapper_717afd68_in;
output	[15:0]	endianswapper_717afd68_out;
assign endianswapper_717afd68_out=endianswapper_717afd68_in;
endmodule



module LL1_L_iunzipFilter2D_endianswapper_2f332b30_(endianswapper_2f332b30_in, endianswapper_2f332b30_out);
input	[15:0]	endianswapper_2f332b30_in;
output	[15:0]	endianswapper_2f332b30_out;
assign endianswapper_2f332b30_out=endianswapper_2f332b30_in;
endmodule



module LL1_L_iunzipFilter2D_stateVar_processedRows(bus_50f9a42f_, bus_2540158d_, bus_029cd39d_, bus_3a105536_, bus_3b123367_, bus_52a23a90_, bus_178131c8_, bus_25bedb97_, bus_1305960f_, bus_7e5a3b31_, bus_6ba6e043_, bus_30eeb15a_, bus_5d02476d_, bus_137b120f_, bus_0d79e859_, bus_406a29e0_, bus_3f13ae55_, bus_707ce562_, bus_7a4ea340_);
input		bus_50f9a42f_;
input		bus_2540158d_;
input		bus_029cd39d_;
input	[15:0]	bus_3a105536_;
input		bus_3b123367_;
input	[15:0]	bus_52a23a90_;
input		bus_178131c8_;
input	[15:0]	bus_25bedb97_;
input		bus_1305960f_;
input	[15:0]	bus_7e5a3b31_;
input		bus_6ba6e043_;
input	[15:0]	bus_30eeb15a_;
input		bus_5d02476d_;
input	[15:0]	bus_137b120f_;
input		bus_0d79e859_;
input	[15:0]	bus_406a29e0_;
input		bus_3f13ae55_;
input	[15:0]	bus_707ce562_;
output	[15:0]	bus_7a4ea340_;
wire	[15:0]	endianswapper_717afd68_out;
reg	[15:0]	stateVar_processedRows_u1=16'h0;
wire	[15:0]	endianswapper_2f332b30_out;
wire		or_7d7f58e7_u0;
wire	[15:0]	mux_21738fda_u0;
LL1_L_iunzipFilter2D_endianswapper_717afd68_ LL1_L_iunzipFilter2D_endianswapper_717afd68__1(.endianswapper_717afd68_in(mux_21738fda_u0), 
  .endianswapper_717afd68_out(endianswapper_717afd68_out));
assign bus_7a4ea340_=endianswapper_2f332b30_out;
always @(posedge bus_50f9a42f_ or posedge bus_2540158d_)
begin
if (bus_2540158d_)
stateVar_processedRows_u1<=16'h0;
else if (or_7d7f58e7_u0)
stateVar_processedRows_u1<=endianswapper_717afd68_out;
end
LL1_L_iunzipFilter2D_endianswapper_2f332b30_ LL1_L_iunzipFilter2D_endianswapper_2f332b30__1(.endianswapper_2f332b30_in(stateVar_processedRows_u1), 
  .endianswapper_2f332b30_out(endianswapper_2f332b30_out));
assign or_7d7f58e7_u0=bus_029cd39d_|bus_3b123367_|bus_178131c8_|bus_1305960f_|bus_6ba6e043_|bus_5d02476d_|bus_0d79e859_|bus_3f13ae55_;
assign mux_21738fda_u0=({16{bus_029cd39d_}}&bus_3a105536_)|({16{bus_3b123367_}}&16'h1)|({16{bus_178131c8_}}&bus_25bedb97_)|({16{bus_1305960f_}}&bus_7e5a3b31_)|({16{bus_6ba6e043_}}&bus_30eeb15a_)|({16{bus_5d02476d_}}&bus_137b120f_)|({16{bus_0d79e859_}}&16'h0)|({16{bus_3f13ae55_}}&16'h0);
endmodule



module LL1_L_iunzipFilter2D_midRightNoConsume2(CLK, RESET, GO, port_79bca4ff_, port_2d1fccd3_, port_79275d09_, port_5fb2661f_, RESULT, RESULT_u691, RESULT_u692, RESULT_u693, RESULT_u694, RESULT_u695, RESULT_u696, RESULT_u697, RESULT_u698, RESULT_u699, RESULT_u700, RESULT_u701, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_79bca4ff_;
input		port_2d1fccd3_;
input		port_79275d09_;
input	[15:0]	port_5fb2661f_;
output		RESULT;
output	[15:0]	RESULT_u691;
output		RESULT_u692;
output	[15:0]	RESULT_u693;
output		RESULT_u694;
output		RESULT_u695;
output		RESULT_u696;
output	[31:0]	RESULT_u697;
output	[2:0]	RESULT_u698;
output	[15:0]	RESULT_u699;
output	[15:0]	RESULT_u700;
output		RESULT_u701;
output		DONE;
wire		and_u1228_u0;
reg		done_cache_u78=1'h0;
wire		or_u327_u0;
wire		or_u328_u0;
reg		done_cache_u79_u0=1'h0;
wire		and_u1233_u0;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_263227c1_instance_RESULT;
wire	[15:0]	add;
wire		not_u237;
wire	[15:0]	simplePinWrite;
wire	[15:0]	simplePinWrite_u194;
wire		simplePinWrite_u195;
reg		reg_24921e83_u0=1'h0;
reg		reg_5e46986b_u0=1'h0;
reg	[15:0]	syncEnable_u59=16'h0;
reg		reg_24921e83_result_delayed_u0=1'h0;
reg		reg_5e46986b_result_delayed_u0=1'h0;
wire		or_u329_u0;
reg		reg_24921e83_result_delayed_result_delayed_u0=1'h0;
assign and_u1228_u0=done_cache_u78&port_79275d09_;
always @(posedge CLK or posedge GO or posedge or_u327_u0)
begin
if (or_u327_u0)
done_cache_u78<=1'h0;
else if (GO)
done_cache_u78<=1'h1;
else done_cache_u78<=done_cache_u78;
end
assign or_u327_u0=and_u1228_u0|RESET;
assign or_u328_u0=and_u1233_u0|RESET;
always @(posedge CLK or posedge reg_5e46986b_result_delayed_u0 or posedge or_u328_u0)
begin
if (or_u328_u0)
done_cache_u79_u0<=1'h0;
else if (reg_5e46986b_result_delayed_u0)
done_cache_u79_u0<=1'h1;
else done_cache_u79_u0<=done_cache_u79_u0;
end
assign and_u1233_u0=done_cache_u79_u0&port_79275d09_;
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_263227c1_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_263227c1_instance(.GO(reg_24921e83_u0), 
  .port_183f8c2f_(syncEnable_u59), .port_7b66f983_(port_5fb2661f_), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_263227c1_instance_RESULT));
assign add=port_79bca4ff_+16'h1;
assign not_u237=!port_2d1fccd3_;
assign simplePinWrite=16'h1&{16{1'h1}};
assign simplePinWrite_u194=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_263227c1_instance_RESULT&{16{reg_24921e83_u0}};
assign simplePinWrite_u195=reg_24921e83_u0&{1{reg_24921e83_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_24921e83_u0<=1'h0;
else reg_24921e83_u0<=reg_5e46986b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5e46986b_u0<=1'h0;
else reg_5e46986b_u0<=GO;
end
always @(posedge CLK)
begin
if (reg_5e46986b_u0)
syncEnable_u59<=port_5fb2661f_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_24921e83_result_delayed_u0<=1'h0;
else reg_24921e83_result_delayed_u0<=reg_24921e83_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5e46986b_result_delayed_u0<=1'h0;
else reg_5e46986b_result_delayed_u0<=reg_5e46986b_u0;
end
assign or_u329_u0=GO|reg_5e46986b_result_delayed_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_24921e83_result_delayed_result_delayed_u0<=1'h0;
else reg_24921e83_result_delayed_result_delayed_u0<=reg_24921e83_result_delayed_u0;
end
assign RESULT=GO;
assign RESULT_u691=add;
assign RESULT_u692=GO;
assign RESULT_u693=16'h0;
assign RESULT_u694=GO;
assign RESULT_u695=not_u237;
assign RESULT_u696=or_u329_u0;
assign RESULT_u697=32'h0;
assign RESULT_u698=3'h1;
assign RESULT_u699=simplePinWrite_u194;
assign RESULT_u700=simplePinWrite;
assign RESULT_u701=simplePinWrite_u195;
assign DONE=reg_24921e83_result_delayed_result_delayed_u0;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_263227c1_(GO, port_183f8c2f_, port_7b66f983_, RESULT);
input		GO;
input	[15:0]	port_183f8c2f_;
input	[15:0]	port_7b66f983_;
output	[15:0]	RESULT;
wire	[15:0]	subtract;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_3511e6d9_instance_RESULT;
assign subtract=port_183f8c2f_-port_7b66f983_;
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_3511e6d9_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_3511e6d9_instance(.GO(GO), 
  .port_5cf61c88_({subtract[15], subtract[15:1]}), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_3511e6d9_instance_RESULT));
assign RESULT=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_3511e6d9_instance_RESULT;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_3511e6d9_(GO, port_5cf61c88_, RESULT);
input		GO;
input	[15:0]	port_5cf61c88_;
output	[15:0]	RESULT;
wire signed	[15:0]	greaterThan_b_signed;
wire signed	[15:0]	greaterThan_a_signed;
wire		greaterThan;
wire		not_u236_u0;
wire		and_u1237_u0;
wire		and_u1238_u0;
wire		and_u1239_u0;
wire	[15:0]	mux_u77;
wire		and_u1240_u0;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_5cf61c88_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign not_u236_u0=~greaterThan;
assign and_u1237_u0=GO&not_u236_u0;
assign and_u1238_u0=GO&greaterThan;
assign and_u1239_u0=and_u1237_u0&GO;
assign mux_u77=(and_u1239_u0)?port_5cf61c88_:16'h0;
assign and_u1240_u0=and_u1238_u0&GO;
assign RESULT=mux_u77;
endmodule



module LL1_L_iunzipFilter2D_endianswapper_0547ae50_(endianswapper_0547ae50_in, endianswapper_0547ae50_out);
input	[31:0]	endianswapper_0547ae50_in;
output	[31:0]	endianswapper_0547ae50_out;
assign endianswapper_0547ae50_out=endianswapper_0547ae50_in;
endmodule



module LL1_L_iunzipFilter2D_endianswapper_4c46d6cc_(endianswapper_4c46d6cc_in, endianswapper_4c46d6cc_out);
input	[31:0]	endianswapper_4c46d6cc_in;
output	[31:0]	endianswapper_4c46d6cc_out;
assign endianswapper_4c46d6cc_out=endianswapper_4c46d6cc_in;
endmodule



module LL1_L_iunzipFilter2D_stateVar_consumed(bus_7424c935_, bus_1123d441_, bus_3f16ffcc_, bus_6227a442_, bus_7b8e9386_, bus_067c086b_, bus_0dde284b_, bus_07d88328_, bus_652ccf5e_, bus_48c0b833_, bus_3323d058_, bus_606ed600_, bus_48687f49_, bus_64ad0da3_, bus_2c867b3c_, bus_7aacda2c_, bus_3c7f9dca_, bus_56028ff8_, bus_4fdd9249_, bus_5dd8910a_, bus_17ac4f32_, bus_2ca297c8_, bus_6b11aeca_, bus_3e36f63b_, bus_4b2a5c22_, bus_55ce97a1_, bus_3d462f24_);
input		bus_7424c935_;
input		bus_1123d441_;
input		bus_3f16ffcc_;
input	[31:0]	bus_6227a442_;
input		bus_7b8e9386_;
input	[31:0]	bus_067c086b_;
input		bus_0dde284b_;
input	[31:0]	bus_07d88328_;
input		bus_652ccf5e_;
input	[31:0]	bus_48c0b833_;
input		bus_3323d058_;
input	[31:0]	bus_606ed600_;
input		bus_48687f49_;
input	[31:0]	bus_64ad0da3_;
input		bus_2c867b3c_;
input	[31:0]	bus_7aacda2c_;
input		bus_3c7f9dca_;
input	[31:0]	bus_56028ff8_;
input		bus_4fdd9249_;
input	[31:0]	bus_5dd8910a_;
input		bus_17ac4f32_;
input	[31:0]	bus_2ca297c8_;
input		bus_6b11aeca_;
input	[31:0]	bus_3e36f63b_;
input		bus_4b2a5c22_;
input	[31:0]	bus_55ce97a1_;
output	[31:0]	bus_3d462f24_;
wire		or_20e6bfa3_u0;
wire	[31:0]	endianswapper_0547ae50_out;
wire	[31:0]	mux_1d9f5947_u0;
reg	[31:0]	stateVar_consumed_u1=32'h0;
wire	[31:0]	endianswapper_4c46d6cc_out;
assign or_20e6bfa3_u0=bus_3f16ffcc_|bus_7b8e9386_|bus_0dde284b_|bus_652ccf5e_|bus_3323d058_|bus_48687f49_|bus_2c867b3c_|bus_3c7f9dca_|bus_4fdd9249_|bus_17ac4f32_|bus_6b11aeca_|bus_4b2a5c22_;
LL1_L_iunzipFilter2D_endianswapper_0547ae50_ LL1_L_iunzipFilter2D_endianswapper_0547ae50__1(.endianswapper_0547ae50_in(mux_1d9f5947_u0), 
  .endianswapper_0547ae50_out(endianswapper_0547ae50_out));
assign mux_1d9f5947_u0=({32{bus_3f16ffcc_}}&bus_6227a442_)|({32{bus_7b8e9386_}}&bus_067c086b_)|({32{bus_0dde284b_}}&bus_07d88328_)|({32{bus_652ccf5e_}}&bus_48c0b833_)|({32{bus_3323d058_}}&bus_606ed600_)|({32{bus_48687f49_}}&bus_64ad0da3_)|({32{bus_2c867b3c_}}&bus_7aacda2c_)|({32{bus_3c7f9dca_}}&bus_56028ff8_)|({32{bus_4fdd9249_}}&bus_5dd8910a_)|({32{bus_17ac4f32_}}&bus_2ca297c8_)|({32{bus_6b11aeca_}}&32'h0)|({32{bus_4b2a5c22_}}&32'h0);
always @(posedge bus_7424c935_ or posedge bus_1123d441_)
begin
if (bus_1123d441_)
stateVar_consumed_u1<=32'h0;
else if (or_20e6bfa3_u0)
stateVar_consumed_u1<=endianswapper_0547ae50_out;
end
LL1_L_iunzipFilter2D_endianswapper_4c46d6cc_ LL1_L_iunzipFilter2D_endianswapper_4c46d6cc__1(.endianswapper_4c46d6cc_in(stateVar_consumed_u1), 
  .endianswapper_4c46d6cc_out(endianswapper_4c46d6cc_out));
assign bus_3d462f24_=endianswapper_4c46d6cc_out;
endmodule



module LL1_L_iunzipFilter2D_endianswapper_543ff5d9_(endianswapper_543ff5d9_in, endianswapper_543ff5d9_out);
input	[2:0]	endianswapper_543ff5d9_in;
output	[2:0]	endianswapper_543ff5d9_out;
assign endianswapper_543ff5d9_out=endianswapper_543ff5d9_in;
endmodule



module LL1_L_iunzipFilter2D_endianswapper_25c43773_(endianswapper_25c43773_in, endianswapper_25c43773_out);
input	[2:0]	endianswapper_25c43773_in;
output	[2:0]	endianswapper_25c43773_out;
assign endianswapper_25c43773_out=endianswapper_25c43773_in;
endmodule



module LL1_L_iunzipFilter2D_stateVar_fsmState_LL1_L_iunzipFilter2D(bus_345dfb8f_, bus_61dd5bb3_, bus_6854f934_, bus_38852323_, bus_5db5252c_);
input		bus_345dfb8f_;
input		bus_61dd5bb3_;
input		bus_6854f934_;
input	[2:0]	bus_38852323_;
output	[2:0]	bus_5db5252c_;
reg	[2:0]	stateVar_fsmState_LL1_L_iunzipFilter2D_u0=3'h0;
wire	[2:0]	endianswapper_543ff5d9_out;
wire	[2:0]	endianswapper_25c43773_out;
always @(posedge bus_345dfb8f_ or posedge bus_61dd5bb3_)
begin
if (bus_61dd5bb3_)
stateVar_fsmState_LL1_L_iunzipFilter2D_u0<=3'h0;
else if (bus_6854f934_)
stateVar_fsmState_LL1_L_iunzipFilter2D_u0<=endianswapper_543ff5d9_out;
end
LL1_L_iunzipFilter2D_endianswapper_543ff5d9_ LL1_L_iunzipFilter2D_endianswapper_543ff5d9__1(.endianswapper_543ff5d9_in(bus_38852323_), 
  .endianswapper_543ff5d9_out(endianswapper_543ff5d9_out));
LL1_L_iunzipFilter2D_endianswapper_25c43773_ LL1_L_iunzipFilter2D_endianswapper_25c43773__1(.endianswapper_25c43773_in(stateVar_fsmState_LL1_L_iunzipFilter2D_u0), 
  .endianswapper_25c43773_out(endianswapper_25c43773_out));
assign bus_5db5252c_=endianswapper_25c43773_out;
endmodule



module LL1_L_iunzipFilter2D_midLeftNoConsume1(CLK, RESET, GO, port_5a8739a4_, port_75d6138f_, port_13e22dd9_, port_78b51d4c_, RESULT, RESULT_u702, RESULT_u703, RESULT_u704, RESULT_u705, RESULT_u706, RESULT_u707, RESULT_u708, RESULT_u709, RESULT_u710, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_5a8739a4_;
input	[15:0]	port_75d6138f_;
input		port_13e22dd9_;
input	[15:0]	port_78b51d4c_;
output		RESULT;
output	[15:0]	RESULT_u702;
output		RESULT_u703;
output	[15:0]	RESULT_u704;
output		RESULT_u705;
output	[31:0]	RESULT_u706;
output	[2:0]	RESULT_u707;
output	[15:0]	RESULT_u708;
output	[15:0]	RESULT_u709;
output		RESULT_u710;
output		DONE;
wire		or_u330_u0;
reg		done_cache_u80=1'h0;
wire		and_u1241_u0;
reg		done_cache_u81_u0=1'h0;
wire		or_u331_u0;
wire		and_u1246_u0;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_69dcaf27_instance_RESULT;
wire	[15:0]	add;
wire		simplePinWrite;
wire	[15:0]	simplePinWrite_u196;
wire	[15:0]	simplePinWrite_u197;
reg		reg_03b0be81_u0=1'h0;
reg		reg_358eeeee_u0=1'h0;
wire		or_u332_u0;
reg		reg_3615c093_u0=1'h0;
reg	[15:0]	syncEnable_u60=16'h0;
reg		reg_0858dc90_u0=1'h0;
reg		reg_03b0be81_result_delayed_u0=1'h0;
assign or_u330_u0=and_u1241_u0|RESET;
always @(posedge CLK or posedge GO or posedge or_u330_u0)
begin
if (or_u330_u0)
done_cache_u80<=1'h0;
else if (GO)
done_cache_u80<=1'h1;
else done_cache_u80<=done_cache_u80;
end
assign and_u1241_u0=done_cache_u80&port_13e22dd9_;
always @(posedge CLK or posedge reg_03b0be81_u0 or posedge or_u331_u0)
begin
if (or_u331_u0)
done_cache_u81_u0<=1'h0;
else if (reg_03b0be81_u0)
done_cache_u81_u0<=1'h1;
else done_cache_u81_u0<=done_cache_u81_u0;
end
assign or_u331_u0=and_u1246_u0|RESET;
assign and_u1246_u0=done_cache_u81_u0&port_13e22dd9_;
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_69dcaf27_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_69dcaf27_instance(.GO(reg_03b0be81_result_delayed_u0), 
  .port_48cd0105_(port_78b51d4c_), .port_047c8d5d_(syncEnable_u60), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_69dcaf27_instance_RESULT));
assign add=port_75d6138f_+16'h1;
assign simplePinWrite=reg_03b0be81_result_delayed_u0&{1{reg_03b0be81_result_delayed_u0}};
assign simplePinWrite_u196=16'h1&{16{1'h1}};
assign simplePinWrite_u197=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_69dcaf27_instance_RESULT&{16{reg_03b0be81_result_delayed_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_03b0be81_u0<=1'h0;
else reg_03b0be81_u0<=reg_0858dc90_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_358eeeee_u0<=1'h0;
else reg_358eeeee_u0<=reg_3615c093_u0;
end
assign or_u332_u0=GO|reg_03b0be81_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3615c093_u0<=1'h0;
else reg_3615c093_u0<=reg_03b0be81_result_delayed_u0;
end
always @(posedge CLK)
begin
if (reg_0858dc90_u0)
syncEnable_u60<=port_78b51d4c_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0858dc90_u0<=1'h0;
else reg_0858dc90_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_03b0be81_result_delayed_u0<=1'h0;
else reg_03b0be81_result_delayed_u0<=reg_03b0be81_u0;
end
assign RESULT=GO;
assign RESULT_u702=16'h0;
assign RESULT_u703=GO;
assign RESULT_u704=add;
assign RESULT_u705=or_u332_u0;
assign RESULT_u706=32'h0;
assign RESULT_u707=3'h1;
assign RESULT_u708=simplePinWrite_u197;
assign RESULT_u709=simplePinWrite_u196;
assign RESULT_u710=simplePinWrite;
assign DONE=reg_358eeeee_u0;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_69dcaf27_(GO, port_48cd0105_, port_047c8d5d_, RESULT);
input		GO;
input	[15:0]	port_48cd0105_;
input	[15:0]	port_047c8d5d_;
output	[15:0]	RESULT;
wire	[16:0]	add;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_7f577b5d_instance_RESULT;
assign add={port_047c8d5d_[15], port_047c8d5d_}+{port_48cd0105_[15], port_48cd0105_};
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_7f577b5d_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_7f577b5d_instance(.GO(GO), 
  .port_37a329a4_({add[16], add[16:2]}), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_7f577b5d_instance_RESULT));
assign RESULT=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_7f577b5d_instance_RESULT;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_7f577b5d_(GO, port_37a329a4_, RESULT);
input		GO;
input	[15:0]	port_37a329a4_;
output	[15:0]	RESULT;
wire		greaterThan;
wire signed	[15:0]	greaterThan_a_signed;
wire signed	[15:0]	greaterThan_b_signed;
wire		not_u238_u0;
wire		and_u1250_u0;
wire		and_u1251_u0;
wire		and_u1252_u0;
wire		and_u1253_u0;
wire	[15:0]	mux_u78;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_37a329a4_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign not_u238_u0=~greaterThan;
assign and_u1250_u0=GO&greaterThan;
assign and_u1251_u0=GO&not_u238_u0;
assign and_u1252_u0=and_u1251_u0&GO;
assign and_u1253_u0=and_u1250_u0&GO;
assign mux_u78=(and_u1252_u0)?port_37a329a4_:16'h0;
assign RESULT=mux_u78;
endmodule



module LL1_L_iunzipFilter2D_midNoConsume2(CLK, RESET, GO, port_0df859e8_, port_3e58b459_, port_14715090_, RESULT, RESULT_u711, RESULT_u712, RESULT_u713, RESULT_u714, RESULT_u715, RESULT_u716, RESULT_u717, RESULT_u718, RESULT_u719, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_0df859e8_;
input		port_3e58b459_;
input	[15:0]	port_14715090_;
output		RESULT;
output	[15:0]	RESULT_u711;
output		RESULT_u712;
output	[15:0]	RESULT_u713;
output		RESULT_u714;
output	[31:0]	RESULT_u715;
output	[2:0]	RESULT_u716;
output	[15:0]	RESULT_u717;
output	[15:0]	RESULT_u718;
output		RESULT_u719;
output		DONE;
reg		done_cache_u82=1'h0;
wire		or_u333_u0;
wire		and_u1256_u0;
wire		or_u334_u0;
wire		and_u1261_u0;
reg		done_cache_u83_u0=1'h0;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_210568e0_instance_RESULT;
wire	[15:0]	add;
wire	[15:0]	simplePinWrite;
wire	[15:0]	simplePinWrite_u198;
wire		simplePinWrite_u199;
reg		reg_3134f12f_u0=1'h0;
reg	[15:0]	syncEnable_u61=16'h0;
reg		reg_505b8c66_u0=1'h0;
reg		reg_5f6fe93d_u0=1'h0;
wire		or_u335_u0;
reg		reg_3134f12f_result_delayed_u0=1'h0;
reg		reg_3134f12f_result_delayed_result_delayed_u0=1'h0;
always @(posedge CLK or posedge GO or posedge or_u333_u0)
begin
if (or_u333_u0)
done_cache_u82<=1'h0;
else if (GO)
done_cache_u82<=1'h1;
else done_cache_u82<=done_cache_u82;
end
assign or_u333_u0=and_u1256_u0|RESET;
assign and_u1256_u0=done_cache_u82&port_3e58b459_;
assign or_u334_u0=and_u1261_u0|RESET;
assign and_u1261_u0=done_cache_u83_u0&port_3e58b459_;
always @(posedge CLK or posedge reg_3134f12f_u0 or posedge or_u334_u0)
begin
if (or_u334_u0)
done_cache_u83_u0<=1'h0;
else if (reg_3134f12f_u0)
done_cache_u83_u0<=1'h1;
else done_cache_u83_u0<=done_cache_u83_u0;
end
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_210568e0_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_210568e0_instance(.GO(reg_3134f12f_result_delayed_u0), 
  .port_27711aa7_(port_14715090_), .port_1d831cf5_(syncEnable_u61), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_210568e0_instance_RESULT));
assign add=port_0df859e8_+16'h1;
assign simplePinWrite=16'h1&{16{1'h1}};
assign simplePinWrite_u198=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_210568e0_instance_RESULT&{16{reg_3134f12f_result_delayed_u0}};
assign simplePinWrite_u199=reg_3134f12f_result_delayed_u0&{1{reg_3134f12f_result_delayed_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3134f12f_u0<=1'h0;
else reg_3134f12f_u0<=reg_505b8c66_u0;
end
always @(posedge CLK)
begin
if (reg_505b8c66_u0)
syncEnable_u61<=port_14715090_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_505b8c66_u0<=1'h0;
else reg_505b8c66_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5f6fe93d_u0<=1'h0;
else reg_5f6fe93d_u0<=reg_3134f12f_result_delayed_result_delayed_u0;
end
assign or_u335_u0=GO|reg_3134f12f_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3134f12f_result_delayed_u0<=1'h0;
else reg_3134f12f_result_delayed_u0<=reg_3134f12f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3134f12f_result_delayed_result_delayed_u0<=1'h0;
else reg_3134f12f_result_delayed_result_delayed_u0<=reg_3134f12f_result_delayed_u0;
end
assign RESULT=GO;
assign RESULT_u711=16'h0;
assign RESULT_u712=GO;
assign RESULT_u713=add;
assign RESULT_u714=or_u335_u0;
assign RESULT_u715=32'h0;
assign RESULT_u716=3'h1;
assign RESULT_u717=simplePinWrite_u198;
assign RESULT_u718=simplePinWrite;
assign RESULT_u719=simplePinWrite_u199;
assign DONE=reg_5f6fe93d_u0;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_210568e0_(GO, port_27711aa7_, port_1d831cf5_, RESULT);
input		GO;
input	[15:0]	port_27711aa7_;
input	[15:0]	port_1d831cf5_;
output	[15:0]	RESULT;
wire	[15:0]	subtract;
wire	[15:0]	LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_563a3424_instance_RESULT;
assign subtract=port_1d831cf5_-port_27711aa7_;
LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_563a3424_ LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_563a3424_instance(.GO(GO), 
  .port_7d7baa57_({subtract[15], subtract[15:1]}), .RESULT(LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_563a3424_instance_RESULT));
assign RESULT=LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_563a3424_instance_RESULT;
endmodule



module LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_LL1_L_iunzipFilter2D_procedure_563a3424_(GO, port_7d7baa57_, RESULT);
input		GO;
input	[15:0]	port_7d7baa57_;
output	[15:0]	RESULT;
wire signed	[15:0]	greaterThan_a_signed;
wire signed	[15:0]	greaterThan_b_signed;
wire		greaterThan;
wire		not_u239_u0;
wire		and_u1265_u0;
wire		and_u1266_u0;
wire		and_u1267_u0;
wire	[15:0]	mux_u79;
wire		and_u1268_u0;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_7d7baa57_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign not_u239_u0=~greaterThan;
assign and_u1265_u0=GO&greaterThan;
assign and_u1266_u0=GO&not_u239_u0;
assign and_u1267_u0=and_u1265_u0&GO;
assign mux_u79=(and_u1267_u0)?16'h0:port_7d7baa57_;
assign and_u1268_u0=and_u1266_u0&GO;
assign RESULT=mux_u79;
endmodule


