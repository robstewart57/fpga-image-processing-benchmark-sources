// __  ___ __ ___  _ __   ___  ___ 
// \ \/ / '__/ _ \| '_ \ / _ \/ __|
//  >  <| | | (_) | | | | (_) \__ \
// /_/\_\_|  \___/|_| |_|\___/|___/
// 
// Xronos synthesizer version
// Run date: Thu 2 Nov 2017 13:58:34 +0000
// 

module LL1_iunzip(Out1_SEND, CLK, In1_COUNT, Out1_DATA, Out1_COUNT, In1_SEND, Out2_ACK, Out2_RDY, In1_DATA, Out1_ACK, RESET, In1_ACK, Out1_RDY, Out2_DATA, Out2_COUNT, Out2_SEND);
output		Out1_SEND;
input		CLK;
wire		streamEndFun1_go;
input	[15:0]	In1_COUNT;
wire		streamFun1_done;
output	[15:0]	Out1_DATA;
output	[15:0]	Out1_COUNT;
input		In1_SEND;
wire		firstNPixels_done;
input		Out2_ACK;
input		Out2_RDY;
wire		streamFun1_go;
wire		streamEndFun1_done;
wire		streamEndFun2_done;
input	[15:0]	In1_DATA;
wire		firstNPixels_go;
input		Out1_ACK;
input		RESET;
output		In1_ACK;
input		Out1_RDY;
wire		streamFun2_done;
wire		streamEndFun2_go;
output	[15:0]	Out2_DATA;
wire		streamFun2_go;
output	[15:0]	Out2_COUNT;
output		Out2_SEND;
wire	[15:0]	streamFun1_u33;
wire		streamFun1_u31;
wire	[31:0]	streamFun1_u28;
wire		streamFun1_u30;
wire		streamFun1_u20;
wire	[2:0]	streamFun1_u23;
wire	[15:0]	streamFun1_u32;
wire		streamFun1_u27;
wire		LL1_iunzip_streamFun1_instance_DONE;
wire		streamFun1;
wire		streamFun1_u18;
wire	[2:0]	streamFun1_u29;
wire	[31:0]	streamFun1_u21;
wire	[31:0]	streamFun1_u19;
wire		streamFun1_u17;
wire		streamFun1_u24;
wire	[31:0]	streamFun1_u25;
wire	[2:0]	streamFun1_u26;
wire	[15:0]	streamFun1_u22;
wire	[31:0]	bus_5e7b48d4_;
wire		bus_1489bd03_;
wire	[2:0]	bus_4f579630_;
wire	[15:0]	bus_3e10c076_;
wire	[31:0]	bus_793d13ac_;
wire		bus_653c2ccc_;
wire	[15:0]	bus_4f4eb58f_;
wire		bus_00a43355_;
wire		bus_2c2b781c_;
wire		bus_69ca0008_;
wire		or_71057e09_u0;
wire		bus_7d0e7909_;
wire		or_05c84b59_u0;
wire		LL1_iunzip_firstNPixels_instance_DONE;
wire	[31:0]	firstNPixels_u11;
wire		firstNPixels_u12;
wire	[31:0]	firstNPixels_u13;
wire	[31:0]	firstNPixels_u19;
wire	[2:0]	firstNPixels_u21;
wire		firstNPixels;
wire	[2:0]	firstNPixels_u14;
wire	[31:0]	firstNPixels_u16;
wire	[2:0]	firstNPixels_u17;
wire		firstNPixels_u15;
wire		firstNPixels_u18;
wire	[15:0]	firstNPixels_u20;
wire		bus_4867c789_;
wire	[15:0]	bus_41de6c42_;
wire		bus_15790327_;
wire	[15:0]	bus_55100efa_;
wire		bus_338070be_;
wire	[15:0]	streamEndFun2_u20;
wire		streamEndFun2;
wire		streamEndFun2_u17;
wire	[2:0]	streamEndFun2_u19;
wire		LL1_iunzip_streamEndFun2_instance_DONE;
wire		streamEndFun2_u21;
wire		streamEndFun2_u25;
wire	[15:0]	streamEndFun2_u22;
wire	[15:0]	streamEndFun2_u24;
wire		streamEndFun2_u14;
wire	[2:0]	streamEndFun2_u16;
wire	[31:0]	streamEndFun2_u18;
wire		streamEndFun2_u13;
wire	[31:0]	streamEndFun2_u15;
wire	[15:0]	streamEndFun2_u23;
wire		bus_251f35c9_;
wire		bus_69d30eb5_;
wire	[15:0]	bus_66064e11_;
wire	[2:0]	bus_1d3e0f48_;
wire		bus_578aeeb2_;
wire		bus_71da01b9_;
wire		bus_17d4c247_;
wire	[15:0]	bus_11305c14_;
wire		bus_4f3b4ae4_;
wire		bus_26f430ba_;
wire	[15:0]	bus_50a40b11_;
wire	[31:0]	bus_2a9ec1c5_;
wire	[15:0]	bus_5c92336e_;
wire		bus_167013f4_;
wire	[15:0]	bus_05a209b3_;
wire	[31:0]	streamFun2_u24;
wire		streamFun2_u20;
wire	[15:0]	streamFun2_u32;
wire		streamFun2;
wire		streamFun2_u17;
wire	[2:0]	streamFun2_u26;
wire	[2:0]	streamFun2_u29;
wire	[31:0]	streamFun2_u21;
wire		streamFun2_u33;
wire		streamFun2_u30;
wire		streamFun2_u27;
wire		streamFun2_u18;
wire	[31:0]	streamFun2_u19;
wire		streamFun2_u23;
wire	[15:0]	streamFun2_u25;
wire		LL1_iunzip_streamFun2_instance_DONE;
wire	[31:0]	streamFun2_u28;
wire	[2:0]	streamFun2_u22;
wire	[15:0]	streamFun2_u31;
wire	[1:0]	bus_7d60e04a_;
wire	[2:0]	bus_306ebd50_;
wire	[15:0]	bus_15657ed6_;
wire	[31:0]	bus_38e2b04c_;
wire		bus_732498ad_;
wire	[15:0]	bus_5a00092e_;
wire		bus_422fb56c_;
wire		bus_7e9b0677_;
wire		bus_26b0e73f_;
wire	[1:0]	bus_3c6b3bea_;
wire	[15:0]	bus_2c07dd11_;
wire	[15:0]	bus_1deedea6_;
wire		bus_0de9df36_;
wire		bus_454c7853_;
wire	[15:0]	or_5ba71816_u0;
wire	[31:0]	bus_22baa6c8_;
wire	[31:0]	bus_072b555f_;
wire		streamEndFun1_u21;
wire	[31:0]	streamEndFun1_u18;
wire	[15:0]	streamEndFun1_u23;
wire	[15:0]	streamEndFun1_u24;
wire	[15:0]	streamEndFun1_u20;
wire	[2:0]	streamEndFun1_u19;
wire		LL1_iunzip_streamEndFun1_instance_DONE;
wire		streamEndFun1_u14;
wire		streamEndFun1_u13;
wire		streamEndFun1_u25;
wire	[31:0]	streamEndFun1_u15;
wire	[2:0]	streamEndFun1_u16;
wire		streamEndFun1_u17;
wire		streamEndFun1;
wire	[15:0]	streamEndFun1_u22;
wire		bus_47c83720_;
wire		bus_35744436_;
wire	[15:0]	bus_3946234b_;
wire		bus_0ace3741_;
wire		bus_6262936b_;
wire	[31:0]	bus_009a4c19_;
wire	[15:0]	bus_69d09001_;
wire	[15:0]	bus_7abd2454_;
wire		bus_23f0e20f_;
wire	[2:0]	bus_1dea0faa_;
wire	[15:0]	bus_1264fa5e_;
wire		bus_7d72a327_;
wire	[15:0]	bus_03be4094_;
wire	[15:0]	or_65ee41bb_u0;
wire		bus_3821ca85_;
wire		or_116b4d36_u0;
wire	[1:0]	scheduler_u111;
wire	[31:0]	scheduler_u115;
wire		scheduler;
wire		scheduler_u119;
wire	[15:0]	scheduler_u122;
wire		scheduler_u125;
wire		scheduler_u126;
wire		scheduler_u116;
wire		scheduler_u114;
wire	[2:0]	scheduler_u123;
wire		scheduler_u128;
wire		scheduler_u112;
wire		LL1_iunzip_scheduler_instance_DONE;
wire	[31:0]	scheduler_u121;
wire		scheduler_u129;
wire		scheduler_u118;
wire	[31:0]	scheduler_u117;
wire		scheduler_u127;
wire	[1:0]	scheduler_u113;
wire		scheduler_u120;
wire		scheduler_u124;
wire	[15:0]	or_18438920_u0;
wire		bus_133bb4de_;
wire		bus_112f1ca0_;
wire	[15:0]	or_380b5f61_u0;
wire		bus_1a0482e7_;
assign Out1_SEND=or_116b4d36_u0;
assign streamEndFun1_go=scheduler_u126;
assign streamFun1_done=bus_3821ca85_;
assign Out1_DATA=or_18438920_u0;
assign Out1_COUNT=or_380b5f61_u0;
assign firstNPixels_done=bus_7d0e7909_;
assign streamFun1_go=scheduler_u125;
assign streamEndFun1_done=bus_112f1ca0_;
assign streamEndFun2_done=bus_133bb4de_;
assign firstNPixels_go=scheduler_u129;
assign In1_ACK=or_71057e09_u0;
assign streamFun2_done=bus_69ca0008_;
assign streamEndFun2_go=scheduler_u127;
assign Out2_DATA=or_65ee41bb_u0;
assign streamFun2_go=scheduler_u128;
assign Out2_COUNT=or_5ba71816_u0;
assign Out2_SEND=or_05c84b59_u0;
LL1_iunzip_streamFun1 LL1_iunzip_streamFun1_instance(.CLK(CLK), .RESET(bus_1a0482e7_), 
  .GO(streamFun1_go), .port_6ca2ba5a_(bus_4867c789_), .port_0abd07fc_(bus_5e7b48d4_), 
  .port_4821e518_(bus_69d30eb5_), .port_57131b69_(bus_69d30eb5_), .port_3cba619a_(bus_5c92336e_), 
  .port_611e8b48_(bus_7d72a327_), .port_093ac5c0_(bus_03be4094_), .port_6b93b5b2_(In1_DATA), 
  .DONE(LL1_iunzip_streamFun1_instance_DONE), .RESULT(streamFun1), .RESULT_u845(streamFun1_u17), 
  .RESULT_u846(streamFun1_u18), .RESULT_u847(streamFun1_u19), .RESULT_u854(streamFun1_u20), 
  .RESULT_u855(streamFun1_u21), .RESULT_u856(streamFun1_u22), .RESULT_u857(streamFun1_u23), 
  .RESULT_u851(streamFun1_u24), .RESULT_u852(streamFun1_u25), .RESULT_u853(streamFun1_u26), 
  .RESULT_u848(streamFun1_u27), .RESULT_u849(streamFun1_u28), .RESULT_u850(streamFun1_u29), 
  .RESULT_u858(streamFun1_u30), .RESULT_u859(streamFun1_u31), .RESULT_u860(streamFun1_u32), 
  .RESULT_u861(streamFun1_u33));
LL1_iunzip_stateVar_consumed LL1_iunzip_stateVar_consumed_1(.bus_40801bcf_(CLK), 
  .bus_4cc978eb_(bus_1a0482e7_), .bus_57fb3572_(firstNPixels), .bus_10ec2e16_(firstNPixels_u11), 
  .bus_63c33e6b_(streamFun1_u18), .bus_2de5c531_(streamFun1_u19), .bus_54819068_(streamFun2_u18), 
  .bus_4dbdf77e_(streamFun2_u19), .bus_5e7b48d4_(bus_5e7b48d4_));
LL1_iunzip_simplememoryreferee_10e4f9e3_ LL1_iunzip_simplememoryreferee_10e4f9e3__1(.bus_4d7cb913_(CLK), 
  .bus_19444fb2_(bus_1a0482e7_), .bus_2b67ea6d_(bus_338070be_), .bus_6066a587_(bus_55100efa_), 
  .bus_3cdb5232_(firstNPixels_u15), .bus_3d51144b_(32'h0), .bus_37d0515c_(3'h1), 
  .bus_4eaf36f8_(scheduler_u120), .bus_4e912bef_(scheduler_u122), .bus_04902313_(scheduler_u121), 
  .bus_2895c6af_(3'h1), .bus_3e10c076_(bus_3e10c076_), .bus_793d13ac_(bus_793d13ac_), 
  .bus_1489bd03_(bus_1489bd03_), .bus_2c2b781c_(bus_2c2b781c_), .bus_4f579630_(bus_4f579630_), 
  .bus_4f4eb58f_(bus_4f4eb58f_), .bus_00a43355_(bus_00a43355_), .bus_653c2ccc_(bus_653c2ccc_));
assign bus_69ca0008_=LL1_iunzip_streamFun2_instance_DONE&{1{LL1_iunzip_streamFun2_instance_DONE}};
assign or_71057e09_u0=streamFun1_u30|streamFun2_u30|scheduler_u124;
assign bus_7d0e7909_=LL1_iunzip_firstNPixels_instance_DONE&{1{LL1_iunzip_firstNPixels_instance_DONE}};
assign or_05c84b59_u0=streamFun2_u33|streamEndFun1_u25|streamEndFun2_u25;
LL1_iunzip_firstNPixels LL1_iunzip_firstNPixels_instance(.CLK(CLK), .RESET(bus_1a0482e7_), 
  .GO(firstNPixels_go), .port_42420f9a_(bus_5e7b48d4_), .port_1b0c101d_(bus_7e9b0677_), 
  .port_735ece5a_(bus_15657ed6_), .port_109251b1_(bus_00a43355_), .port_2f0a27cf_(bus_4f4eb58f_), 
  .port_463aad8f_(bus_26f430ba_), .DONE(LL1_iunzip_firstNPixels_instance_DONE), 
  .RESULT(firstNPixels), .RESULT_u862(firstNPixels_u11), .RESULT_u863(firstNPixels_u12), 
  .RESULT_u864(firstNPixels_u13), .RESULT_u865(firstNPixels_u14), .RESULT_u866(firstNPixels_u15), 
  .RESULT_u867(firstNPixels_u16), .RESULT_u868(firstNPixels_u17), .RESULT_u869(firstNPixels_u18), 
  .RESULT_u870(firstNPixels_u19), .RESULT_u871(firstNPixels_u20), .RESULT_u872(firstNPixels_u21));
LL1_iunzip_stateVar_midPoint LL1_iunzip_stateVar_midPoint_1(.bus_728f42fb_(CLK), 
  .bus_20ca5157_(bus_1a0482e7_), .bus_036aef22_(streamFun1), .bus_794845ef_(1'h0), 
  .bus_36d74eeb_(streamFun2), .bus_51440103_(1'h0), .bus_3a6cc6f4_(streamEndFun1), 
  .bus_63d56c2a_(1'h0), .bus_0a115faf_(streamEndFun2), .bus_110dbdeb_(1'h0), .bus_4867c789_(bus_4867c789_));
LL1_iunzip_structuralmemory_199cf187_ LL1_iunzip_structuralmemory_199cf187__1(.CLK_u4(CLK), 
  .bus_5451230e_(bus_1a0482e7_), .bus_71688263_(32'h1), .bus_7304c986_(3'h1), .bus_3e8fafd7_(bus_732498ad_), 
  .bus_4e7a128c_(bus_793d13ac_), .bus_069ded29_(3'h1), .bus_016e515e_(bus_2c2b781c_), 
  .bus_261f279e_(bus_1489bd03_), .bus_2558522d_(bus_3e10c076_), .bus_41de6c42_(bus_41de6c42_), 
  .bus_15790327_(bus_15790327_), .bus_55100efa_(bus_55100efa_), .bus_338070be_(bus_338070be_));
LL1_iunzip_streamEndFun2 LL1_iunzip_streamEndFun2_instance(.CLK(CLK), .RESET(bus_1a0482e7_), 
  .GO(streamEndFun2_go), .port_3f8bef0c_(bus_4867c789_), .port_59348860_(bus_71da01b9_), 
  .port_38c4f7d8_(bus_66064e11_), .port_3c3e7cb8_(bus_0ace3741_), .port_74b582d8_(bus_7abd2454_), 
  .DONE(LL1_iunzip_streamEndFun2_instance_DONE), .RESULT(streamEndFun2), .RESULT_u873(streamEndFun2_u13), 
  .RESULT_u877(streamEndFun2_u14), .RESULT_u878(streamEndFun2_u15), .RESULT_u879(streamEndFun2_u16), 
  .RESULT_u874(streamEndFun2_u17), .RESULT_u875(streamEndFun2_u18), .RESULT_u876(streamEndFun2_u19), 
  .RESULT_u880(streamEndFun2_u20), .RESULT_u881(streamEndFun2_u21), .RESULT_u882(streamEndFun2_u22), 
  .RESULT_u883(streamEndFun2_u23), .RESULT_u884(streamEndFun2_u24), .RESULT_u885(streamEndFun2_u25));
LL1_iunzip_Kicker_26 LL1_iunzip_Kicker_26_1(.CLK(CLK), .RESET(bus_1a0482e7_), .bus_251f35c9_(bus_251f35c9_));
LL1_iunzip_simplememoryreferee_52a82a09_ LL1_iunzip_simplememoryreferee_52a82a09__1(.bus_2453e19e_(CLK), 
  .bus_1b3c311c_(bus_1a0482e7_), .bus_06bb3bca_(bus_454c7853_), .bus_7f823762_(bus_2c07dd11_), 
  .bus_33f699d7_(firstNPixels_u18), .bus_0e87d9ae_(firstNPixels_u20), .bus_51e962ad_({31'b0, firstNPixels_u19[0]}), 
  .bus_43cb9bbb_(3'h1), .bus_5be4b948_(streamFun1_u24), .bus_238bf419_(streamFun1_u20), 
  .bus_7bd172a7_(streamFun1_u22), .bus_0319de32_(streamFun1_u21), .bus_60a35d69_(3'h1), 
  .bus_7475072e_(streamFun2_u27), .bus_7cd5d094_(streamFun2_u23), .bus_2e6c9d65_(streamFun2_u25), 
  .bus_735b4165_(streamFun2_u24), .bus_2da416ce_(3'h1), .bus_455d1534_(streamEndFun1_u14), 
  .bus_5347953e_(streamEndFun1_u15), .bus_1ebd7ee4_(3'h1), .bus_707f0c59_(streamEndFun2_u14), 
  .bus_1ec36984_(streamEndFun2_u15), .bus_5239f197_(3'h1), .bus_11305c14_(bus_11305c14_), 
  .bus_2a9ec1c5_(bus_2a9ec1c5_), .bus_578aeeb2_(bus_578aeeb2_), .bus_17d4c247_(bus_17d4c247_), 
  .bus_1d3e0f48_(bus_1d3e0f48_), .bus_26f430ba_(bus_26f430ba_), .bus_5c92336e_(bus_5c92336e_), 
  .bus_69d30eb5_(bus_69d30eb5_), .bus_05a209b3_(bus_05a209b3_), .bus_4f3b4ae4_(bus_4f3b4ae4_), 
  .bus_50a40b11_(bus_50a40b11_), .bus_167013f4_(bus_167013f4_), .bus_66064e11_(bus_66064e11_), 
  .bus_71da01b9_(bus_71da01b9_));
LL1_iunzip_streamFun2 LL1_iunzip_streamFun2_instance(.CLK(CLK), .RESET(bus_1a0482e7_), 
  .GO(streamFun2_go), .port_4b4b2561_(bus_4867c789_), .port_5a2a759b_(bus_5e7b48d4_), 
  .port_741f83f2_(bus_47c83720_), .port_3d5a0933_(bus_3946234b_), .port_15d252f1_(bus_4f3b4ae4_), 
  .port_6091a1b3_(bus_4f3b4ae4_), .port_3f9a965b_(bus_05a209b3_), .port_189d0bed_(In1_DATA), 
  .DONE(LL1_iunzip_streamFun2_instance_DONE), .RESULT(streamFun2), .RESULT_u886(streamFun2_u17), 
  .RESULT_u887(streamFun2_u18), .RESULT_u888(streamFun2_u19), .RESULT_u889(streamFun2_u20), 
  .RESULT_u890(streamFun2_u21), .RESULT_u891(streamFun2_u22), .RESULT_u895(streamFun2_u23), 
  .RESULT_u896(streamFun2_u24), .RESULT_u897(streamFun2_u25), .RESULT_u898(streamFun2_u26), 
  .RESULT_u892(streamFun2_u27), .RESULT_u893(streamFun2_u28), .RESULT_u894(streamFun2_u29), 
  .RESULT_u899(streamFun2_u30), .RESULT_u900(streamFun2_u31), .RESULT_u901(streamFun2_u32), 
  .RESULT_u902(streamFun2_u33));
LL1_iunzip_stateVar_fsmOldState_LL1_iunzip LL1_iunzip_stateVar_fsmOldState_LL1_iunzip_1(.bus_20ec10f4_(CLK), 
  .bus_09f76d0f_(bus_1a0482e7_), .bus_7508f03a_(scheduler), .bus_078eb971_(scheduler_u111), 
  .bus_7d60e04a_(bus_7d60e04a_));
LL1_iunzip_simplememoryreferee_7e53def4_ LL1_iunzip_simplememoryreferee_7e53def4__1(.bus_5e9a9b98_(CLK), 
  .bus_0b4a27a7_(bus_1a0482e7_), .bus_6ceb0c3b_(bus_15790327_), .bus_3ec3c7a3_(bus_41de6c42_), 
  .bus_50a4ddaf_(firstNPixels_u12), .bus_04a67922_(32'h1), .bus_40e70fc3_(3'h1), 
  .bus_5a00092e_(bus_5a00092e_), .bus_38e2b04c_(bus_38e2b04c_), .bus_422fb56c_(bus_422fb56c_), 
  .bus_732498ad_(bus_732498ad_), .bus_306ebd50_(bus_306ebd50_), .bus_15657ed6_(bus_15657ed6_), 
  .bus_7e9b0677_(bus_7e9b0677_));
LL1_iunzip_stateVar_In1PortEnable LL1_iunzip_stateVar_In1PortEnable_1(.bus_482b48c2_(CLK), 
  .bus_414ca731_(bus_1a0482e7_), .bus_27b57e02_(scheduler_u118), .bus_119b13c9_(scheduler_u119), 
  .bus_26b0e73f_(bus_26b0e73f_));
LL1_iunzip_stateVar_fsmState_LL1_iunzip LL1_iunzip_stateVar_fsmState_LL1_iunzip_1(.bus_781a7383_(CLK), 
  .bus_11069aeb_(bus_1a0482e7_), .bus_2457321f_(scheduler_u112), .bus_2a0ed9bb_(scheduler_u113), 
  .bus_3c6b3bea_(bus_3c6b3bea_));
LL1_iunzip_structuralmemory_65c92979_ LL1_iunzip_structuralmemory_65c92979__1(.CLK_u5(CLK), 
  .bus_1dee1645_(bus_1a0482e7_), .bus_36216417_(bus_009a4c19_), .bus_06d309bc_(3'h1), 
  .bus_6296f247_(bus_35744436_), .bus_083d81f6_(bus_2a9ec1c5_), .bus_3786b3c5_(3'h1), 
  .bus_0f87e737_(bus_17d4c247_), .bus_7a6a921b_(bus_578aeeb2_), .bus_2c10caec_(bus_11305c14_), 
  .bus_1deedea6_(bus_1deedea6_), .bus_0de9df36_(bus_0de9df36_), .bus_2c07dd11_(bus_2c07dd11_), 
  .bus_454c7853_(bus_454c7853_));
assign or_5ba71816_u0=streamFun2_u32|streamEndFun1_u24|streamEndFun2_u24;
LL1_iunzip_stateVar_In1TokenIndex LL1_iunzip_stateVar_In1TokenIndex_1(.bus_028bcee6_(CLK), 
  .bus_3ce31b6e_(bus_1a0482e7_), .bus_3da9e3d5_(scheduler_u114), .bus_4515a94c_(scheduler_u115), 
  .bus_22baa6c8_(bus_22baa6c8_));
LL1_iunzip_stateVar_In1MaxTokenIndex LL1_iunzip_stateVar_In1MaxTokenIndex_1(.bus_21b70cb9_(CLK), 
  .bus_0a95df40_(bus_1a0482e7_), .bus_68994182_(scheduler_u116), .bus_5519f449_({scheduler_u117[31:2], 1'b0, scheduler_u117[0]}), 
  .bus_072b555f_(bus_072b555f_));
LL1_iunzip_streamEndFun1 LL1_iunzip_streamEndFun1_instance(.CLK(CLK), .RESET(bus_1a0482e7_), 
  .GO(streamEndFun1_go), .port_3b9b03c5_(bus_4867c789_), .port_2d39d825_(bus_167013f4_), 
  .port_768c8415_(bus_50a40b11_), .port_53886836_(bus_23f0e20f_), .port_63c1f3c3_(bus_69d09001_), 
  .DONE(LL1_iunzip_streamEndFun1_instance_DONE), .RESULT(streamEndFun1), .RESULT_u903(streamEndFun1_u13), 
  .RESULT_u907(streamEndFun1_u14), .RESULT_u908(streamEndFun1_u15), .RESULT_u909(streamEndFun1_u16), 
  .RESULT_u904(streamEndFun1_u17), .RESULT_u905(streamEndFun1_u18), .RESULT_u906(streamEndFun1_u19), 
  .RESULT_u910(streamEndFun1_u20), .RESULT_u911(streamEndFun1_u21), .RESULT_u912(streamEndFun1_u22), 
  .RESULT_u913(streamEndFun1_u23), .RESULT_u914(streamEndFun1_u24), .RESULT_u915(streamEndFun1_u25));
LL1_iunzip_simplememoryreferee_1c6f7bbb_ LL1_iunzip_simplememoryreferee_1c6f7bbb__1(.bus_46f786f5_(CLK), 
  .bus_3dd26b70_(bus_1a0482e7_), .bus_31d8e4db_(bus_0de9df36_), .bus_7604351c_(bus_1deedea6_), 
  .bus_4e6481ad_(streamFun1_u27), .bus_6be83458_(streamFun1_u28), .bus_2164d186_(3'h1), 
  .bus_51c5d9cf_(streamFun2_u20), .bus_010f6c42_(streamFun2_u21), .bus_675cdef9_(3'h1), 
  .bus_6f27dbf2_(streamEndFun1_u17), .bus_7943488e_(streamEndFun1_u18), .bus_5c945c19_(3'h1), 
  .bus_5ef9551e_(streamEndFun2_u17), .bus_358645e2_(streamEndFun2_u18), .bus_361af4ce_(3'h1), 
  .bus_1264fa5e_(bus_1264fa5e_), .bus_009a4c19_(bus_009a4c19_), .bus_6262936b_(bus_6262936b_), 
  .bus_35744436_(bus_35744436_), .bus_1dea0faa_(bus_1dea0faa_), .bus_03be4094_(bus_03be4094_), 
  .bus_7d72a327_(bus_7d72a327_), .bus_3946234b_(bus_3946234b_), .bus_47c83720_(bus_47c83720_), 
  .bus_69d09001_(bus_69d09001_), .bus_23f0e20f_(bus_23f0e20f_), .bus_7abd2454_(bus_7abd2454_), 
  .bus_0ace3741_(bus_0ace3741_));
assign or_65ee41bb_u0=streamFun2_u31|streamEndFun1_u20|streamEndFun2_u20;
assign bus_3821ca85_=LL1_iunzip_streamFun1_instance_DONE&{1{LL1_iunzip_streamFun1_instance_DONE}};
assign or_116b4d36_u0=streamFun1_u31|streamEndFun1_u21|streamEndFun2_u21;
LL1_iunzip_scheduler LL1_iunzip_scheduler_instance(.CLK(CLK), .RESET(bus_1a0482e7_), 
  .GO(bus_251f35c9_), .port_42a101cc_(bus_7d60e04a_), .port_711c21e7_(bus_3c6b3bea_), 
  .port_305d8ba1_(bus_22baa6c8_), .port_71394b75_(bus_072b555f_), .port_764c2d23_(bus_5e7b48d4_), 
  .port_1d25b47a_(bus_653c2ccc_), .port_21a66f1f_(In1_SEND), .port_7fc5701f_(firstNPixels_done), 
  .port_22a38371_(Out1_RDY), .port_31572f8d_(Out2_RDY), .port_411771b7_(streamFun1_done), 
  .port_1b55da6d_(streamFun2_done), .port_10bcdaa8_(streamEndFun1_done), .port_0379561c_(streamEndFun2_done), 
  .port_7b10a081_(In1_DATA), .DONE(LL1_iunzip_scheduler_instance_DONE), .RESULT(scheduler), 
  .RESULT_u916(scheduler_u111), .RESULT_u917(scheduler_u112), .RESULT_u918(scheduler_u113), 
  .RESULT_u919(scheduler_u114), .RESULT_u920(scheduler_u115), .RESULT_u921(scheduler_u116), 
  .RESULT_u922(scheduler_u117), .RESULT_u923(scheduler_u118), .RESULT_u924(scheduler_u119), 
  .RESULT_u925(scheduler_u120), .RESULT_u926(scheduler_u121), .RESULT_u927(scheduler_u122), 
  .RESULT_u928(scheduler_u123), .RESULT_u929(scheduler_u124), .RESULT_u930(scheduler_u125), 
  .RESULT_u931(scheduler_u126), .RESULT_u932(scheduler_u127), .RESULT_u933(scheduler_u128), 
  .RESULT_u934(scheduler_u129));
assign or_18438920_u0=streamFun1_u32|streamEndFun1_u22|streamEndFun2_u22;
assign bus_133bb4de_=LL1_iunzip_streamEndFun2_instance_DONE&{1{LL1_iunzip_streamEndFun2_instance_DONE}};
assign bus_112f1ca0_=LL1_iunzip_streamEndFun1_instance_DONE&{1{LL1_iunzip_streamEndFun1_instance_DONE}};
assign or_380b5f61_u0=streamFun1_u33|streamEndFun1_u23|streamEndFun2_u23;
LL1_iunzip_globalreset_physical_7bb59c58_ LL1_iunzip_globalreset_physical_7bb59c58__1(.bus_0bf03daf_(CLK), 
  .bus_7876706a_(RESET), .bus_1a0482e7_(bus_1a0482e7_));
endmodule



module LL1_iunzip_streamFun1(CLK, RESET, GO, port_6ca2ba5a_, port_0abd07fc_, port_611e8b48_, port_093ac5c0_, port_57131b69_, port_3cba619a_, port_4821e518_, port_6b93b5b2_, RESULT, RESULT_u845, RESULT_u846, RESULT_u847, RESULT_u848, RESULT_u849, RESULT_u850, RESULT_u851, RESULT_u852, RESULT_u853, RESULT_u854, RESULT_u855, RESULT_u856, RESULT_u857, RESULT_u858, RESULT_u859, RESULT_u860, RESULT_u861, DONE);
input		CLK;
input		RESET;
input		GO;
input		port_6ca2ba5a_;
input	[31:0]	port_0abd07fc_;
input		port_611e8b48_;
input	[15:0]	port_093ac5c0_;
input		port_57131b69_;
input	[15:0]	port_3cba619a_;
input		port_4821e518_;
input	[15:0]	port_6b93b5b2_;
output		RESULT;
output		RESULT_u845;
output		RESULT_u846;
output	[31:0]	RESULT_u847;
output		RESULT_u848;
output	[31:0]	RESULT_u849;
output	[2:0]	RESULT_u850;
output		RESULT_u851;
output	[31:0]	RESULT_u852;
output	[2:0]	RESULT_u853;
output		RESULT_u854;
output	[31:0]	RESULT_u855;
output	[15:0]	RESULT_u856;
output	[2:0]	RESULT_u857;
output		RESULT_u858;
output		RESULT_u859;
output	[15:0]	RESULT_u860;
output	[15:0]	RESULT_u861;
output		DONE;
wire		simplePinWrite;
wire		or_u387_u0;
reg		reg_2bb11662_u0=1'h0;
wire		and_u1447_u0;
wire	[31:0]	add;
wire		and_u1448_u0;
wire	[8:0]	subtract;
wire		greaterThanEqualTo;
wire signed	[8:0]	greaterThanEqualTo_b_signed;
wire signed	[8:0]	greaterThanEqualTo_a_signed;
wire		and_u1449_u0;
wire		not_u280_u0;
wire		and_u1450_u0;
wire	[8:0]	subtract_u6;
wire		and_u1451_u0;
wire	[8:0]	mux_u113;
wire		and_u1452_u0;
wire	[31:0]	add_u37;
wire		and_u1453_u0;
wire		and_u1455_u0;
wire	[16:0]	add_u38;
wire	[15:0]	subtract_u7;
wire	[31:0]	add_u39;
wire	[15:0]	simplePinWrite_u242;
wire	[15:0]	simplePinWrite_u243;
wire		simplePinWrite_u244;
reg	[31:0]	syncEnable_u101=32'h0;
reg	[15:0]	syncEnable_u102_u0=16'h0;
reg	[15:0]	syncEnable_u103_u0=16'h0;
reg		reg_65099414_u0=1'h0;
reg		reg_6e8f8aab_u0=1'h0;
wire	[31:0]	mux_u114_u0;
wire	[31:0]	mux_u115_u0;
wire		or_u388_u0;
reg	[31:0]	syncEnable_u104_u0=32'h0;
reg		reg_65099414_result_delayed_u0=1'h0;
reg	[15:0]	syncEnable_u105_u0=16'h0;
assign simplePinWrite=GO&{1{GO}};
assign or_u387_u0=and_u1447_u0|RESET;
always @(posedge CLK or posedge reg_65099414_u0 or posedge or_u387_u0)
begin
if (or_u387_u0)
reg_2bb11662_u0<=1'h0;
else if (reg_65099414_u0)
reg_2bb11662_u0<=1'h1;
else reg_2bb11662_u0<=reg_2bb11662_u0;
end
assign and_u1447_u0=reg_2bb11662_u0&port_4821e518_;
assign add={31'b0, port_6ca2ba5a_}+32'h0;
assign and_u1448_u0=reg_65099414_result_delayed_u0&port_611e8b48_;
assign subtract={8'b0, port_6ca2ba5a_}-9'h1;
assign greaterThanEqualTo_a_signed={subtract[2], subtract[2], subtract[2], subtract[2], subtract[2], subtract[2], subtract[2:0]};
assign greaterThanEqualTo_b_signed=9'h0;
assign greaterThanEqualTo=greaterThanEqualTo_a_signed>=greaterThanEqualTo_b_signed;
assign and_u1449_u0=GO&not_u280_u0;
assign not_u280_u0=~greaterThanEqualTo;
assign and_u1450_u0=GO&greaterThanEqualTo;
assign subtract_u6={8'b0, port_6ca2ba5a_}-9'h1;
assign and_u1451_u0=and_u1450_u0&GO;
assign mux_u113=(and_u1451_u0)?{subtract_u6[2], subtract_u6[2], subtract_u6[2], subtract_u6[2], subtract_u6[2], subtract_u6[2], subtract_u6[2:0]}:9'h2;
assign and_u1452_u0=and_u1449_u0&GO;
assign add_u37={mux_u113[2], mux_u113[2], mux_u113[2], mux_u113[2], mux_u113[2], mux_u113[2], mux_u113[2], mux_u113[2], mux_u113[2], mux_u113[2], mux_u113[2], mux_u113[2], mux_u113[2], mux_u113[2], mux_u113[2], mux_u113[2], mux_u113[2], mux_u113[2], mux_u113[2], mux_u113[2], mux_u113[2], mux_u113[2], mux_u113[2], mux_u113[2], mux_u113[2], mux_u113[2], mux_u113[2], mux_u113[2], mux_u113[2], mux_u113[2:0]}+32'h0;
assign and_u1453_u0=reg_65099414_result_delayed_u0&port_4821e518_;
assign and_u1455_u0=reg_6e8f8aab_u0&port_611e8b48_;
assign add_u38={syncEnable_u105_u0[15], syncEnable_u105_u0}+{port_093ac5c0_[15], port_093ac5c0_};
assign subtract_u7=syncEnable_u102_u0-add_u38[16:1];
assign add_u39=port_0abd07fc_+32'h1;
assign simplePinWrite_u242=subtract_u7&{16{reg_6e8f8aab_u0}};
assign simplePinWrite_u243=16'h1&{16{1'h1}};
assign simplePinWrite_u244=reg_6e8f8aab_u0&{1{reg_6e8f8aab_u0}};
always @(posedge CLK)
begin
if (GO)
syncEnable_u101<={add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2:0]};
end
always @(posedge CLK)
begin
if (reg_65099414_result_delayed_u0)
syncEnable_u102_u0<=port_093ac5c0_;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u103_u0<=port_6b93b5b2_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_65099414_u0<=1'h0;
else reg_65099414_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6e8f8aab_u0<=1'h0;
else reg_6e8f8aab_u0<=reg_65099414_result_delayed_u0;
end
assign mux_u114_u0=(reg_65099414_u0)?32'h0:syncEnable_u104_u0;
assign mux_u115_u0=(reg_65099414_result_delayed_u0)?syncEnable_u101:32'h0;
assign or_u388_u0=reg_65099414_result_delayed_u0|reg_6e8f8aab_u0;
always @(posedge CLK)
begin
if (GO)
syncEnable_u104_u0<=add_u37;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_65099414_result_delayed_u0<=1'h0;
else reg_65099414_result_delayed_u0<=reg_65099414_u0;
end
always @(posedge CLK)
begin
if (reg_65099414_result_delayed_u0)
syncEnable_u105_u0<=port_3cba619a_;
end
assign RESULT=GO;
assign RESULT_u845=1'h0;
assign RESULT_u846=GO;
assign RESULT_u847=add_u39;
assign RESULT_u848=or_u388_u0;
assign RESULT_u849=mux_u115_u0;
assign RESULT_u850=3'h1;
assign RESULT_u851=reg_65099414_result_delayed_u0;
assign RESULT_u852=mux_u114_u0;
assign RESULT_u853=3'h1;
assign RESULT_u854=reg_65099414_u0;
assign RESULT_u855=mux_u114_u0;
assign RESULT_u856=syncEnable_u103_u0;
assign RESULT_u857=3'h1;
assign RESULT_u858=simplePinWrite;
assign RESULT_u859=simplePinWrite_u244;
assign RESULT_u860=simplePinWrite_u242;
assign RESULT_u861=simplePinWrite_u243;
assign DONE=reg_6e8f8aab_u0;
endmodule



module LL1_iunzip_endianswapper_06af5a46_(endianswapper_06af5a46_in, endianswapper_06af5a46_out);
input	[31:0]	endianswapper_06af5a46_in;
output	[31:0]	endianswapper_06af5a46_out;
assign endianswapper_06af5a46_out=endianswapper_06af5a46_in;
endmodule



module LL1_iunzip_endianswapper_1a51c85e_(endianswapper_1a51c85e_in, endianswapper_1a51c85e_out);
input	[31:0]	endianswapper_1a51c85e_in;
output	[31:0]	endianswapper_1a51c85e_out;
assign endianswapper_1a51c85e_out=endianswapper_1a51c85e_in;
endmodule



module LL1_iunzip_stateVar_consumed(bus_40801bcf_, bus_4cc978eb_, bus_57fb3572_, bus_10ec2e16_, bus_63c33e6b_, bus_2de5c531_, bus_54819068_, bus_4dbdf77e_, bus_5e7b48d4_);
input		bus_40801bcf_;
input		bus_4cc978eb_;
input		bus_57fb3572_;
input	[31:0]	bus_10ec2e16_;
input		bus_63c33e6b_;
input	[31:0]	bus_2de5c531_;
input		bus_54819068_;
input	[31:0]	bus_4dbdf77e_;
output	[31:0]	bus_5e7b48d4_;
wire		or_400b7268_u0;
reg	[31:0]	stateVar_consumed_u3=32'h0;
wire	[31:0]	mux_11d192e5_u0;
wire	[31:0]	endianswapper_06af5a46_out;
wire	[31:0]	endianswapper_1a51c85e_out;
assign or_400b7268_u0=bus_57fb3572_|bus_63c33e6b_|bus_54819068_;
always @(posedge bus_40801bcf_ or posedge bus_4cc978eb_)
begin
if (bus_4cc978eb_)
stateVar_consumed_u3<=32'h0;
else if (or_400b7268_u0)
stateVar_consumed_u3<=endianswapper_1a51c85e_out;
end
assign mux_11d192e5_u0=({32{bus_57fb3572_}}&bus_10ec2e16_)|({32{bus_63c33e6b_}}&bus_2de5c531_)|({32{bus_54819068_}}&bus_4dbdf77e_);
LL1_iunzip_endianswapper_06af5a46_ LL1_iunzip_endianswapper_06af5a46__1(.endianswapper_06af5a46_in(stateVar_consumed_u3), 
  .endianswapper_06af5a46_out(endianswapper_06af5a46_out));
assign bus_5e7b48d4_=endianswapper_06af5a46_out;
LL1_iunzip_endianswapper_1a51c85e_ LL1_iunzip_endianswapper_1a51c85e__1(.endianswapper_1a51c85e_in(mux_11d192e5_u0), 
  .endianswapper_1a51c85e_out(endianswapper_1a51c85e_out));
endmodule



module LL1_iunzip_simplememoryreferee_10e4f9e3_(bus_4d7cb913_, bus_19444fb2_, bus_2b67ea6d_, bus_6066a587_, bus_3cdb5232_, bus_3d51144b_, bus_37d0515c_, bus_4eaf36f8_, bus_4e912bef_, bus_04902313_, bus_2895c6af_, bus_3e10c076_, bus_793d13ac_, bus_1489bd03_, bus_2c2b781c_, bus_4f579630_, bus_4f4eb58f_, bus_00a43355_, bus_653c2ccc_);
input		bus_4d7cb913_;
input		bus_19444fb2_;
input		bus_2b67ea6d_;
input	[15:0]	bus_6066a587_;
input		bus_3cdb5232_;
input	[31:0]	bus_3d51144b_;
input	[2:0]	bus_37d0515c_;
input		bus_4eaf36f8_;
input	[15:0]	bus_4e912bef_;
input	[31:0]	bus_04902313_;
input	[2:0]	bus_2895c6af_;
output	[15:0]	bus_3e10c076_;
output	[31:0]	bus_793d13ac_;
output		bus_1489bd03_;
output		bus_2c2b781c_;
output	[2:0]	bus_4f579630_;
output	[15:0]	bus_4f4eb58f_;
output		bus_00a43355_;
output		bus_653c2ccc_;
wire		and_71cfc94c_u0;
reg		done_qual_u53=1'h0;
reg		done_qual_u54_u0=1'h0;
wire	[31:0]	mux_0ae111b1_u0;
wire		or_3c0d2e7d_u0;
wire	[15:0]	mux_6d1772e3_u0;
wire		and_641cbb24_u0;
wire		not_2de3519a_u0;
wire		not_254d91b1_u0;
wire		or_57f90cc4_u0;
wire		or_1551232f_u0;
assign and_71cfc94c_u0=or_1551232f_u0&bus_2b67ea6d_;
always @(posedge bus_4d7cb913_)
begin
if (bus_19444fb2_)
done_qual_u53<=1'h0;
else done_qual_u53<=bus_3cdb5232_;
end
always @(posedge bus_4d7cb913_)
begin
if (bus_19444fb2_)
done_qual_u54_u0<=1'h0;
else done_qual_u54_u0<=bus_4eaf36f8_;
end
assign mux_0ae111b1_u0=(bus_3cdb5232_)?32'h0:bus_04902313_;
assign or_3c0d2e7d_u0=bus_4eaf36f8_|done_qual_u54_u0;
assign mux_6d1772e3_u0=({16{bus_4eaf36f8_}}&bus_4e912bef_);
assign bus_3e10c076_=mux_6d1772e3_u0;
assign bus_793d13ac_=mux_0ae111b1_u0;
assign bus_1489bd03_=bus_4eaf36f8_;
assign bus_2c2b781c_=or_57f90cc4_u0;
assign bus_4f579630_=3'h1;
assign bus_4f4eb58f_=bus_6066a587_;
assign bus_00a43355_=and_71cfc94c_u0;
assign bus_653c2ccc_=and_641cbb24_u0;
assign and_641cbb24_u0=or_3c0d2e7d_u0&bus_2b67ea6d_;
assign not_2de3519a_u0=~bus_2b67ea6d_;
assign not_254d91b1_u0=~bus_2b67ea6d_;
assign or_57f90cc4_u0=bus_3cdb5232_|bus_4eaf36f8_;
assign or_1551232f_u0=bus_3cdb5232_|done_qual_u53;
endmodule



module LL1_iunzip_firstNPixels(CLK, RESET, GO, port_42420f9a_, port_1b0c101d_, port_735ece5a_, port_109251b1_, port_2f0a27cf_, port_463aad8f_, RESULT, RESULT_u862, RESULT_u863, RESULT_u864, RESULT_u865, RESULT_u866, RESULT_u867, RESULT_u868, RESULT_u869, RESULT_u870, RESULT_u871, RESULT_u872, DONE);
input		CLK;
input		RESET;
input		GO;
input	[31:0]	port_42420f9a_;
input		port_1b0c101d_;
input	[15:0]	port_735ece5a_;
input		port_109251b1_;
input	[15:0]	port_2f0a27cf_;
input		port_463aad8f_;
output		RESULT;
output	[31:0]	RESULT_u862;
output		RESULT_u863;
output	[31:0]	RESULT_u864;
output	[2:0]	RESULT_u865;
output		RESULT_u866;
output	[31:0]	RESULT_u867;
output	[2:0]	RESULT_u868;
output		RESULT_u869;
output	[31:0]	RESULT_u870;
output	[15:0]	RESULT_u871;
output	[2:0]	RESULT_u872;
output		DONE;
wire		and_u1457_u0;
wire		and_u1458_u0;
wire	[31:0]	add;
wire		and_u1459_u0;
wire		or_u389_u0;
reg		reg_712a5581_u0=1'h0;
wire		or_u390_u0;
wire		and_u1460_u0;
reg		reg_19ab1be5_u0=1'h0;
reg	[15:0]	syncEnable_u106=16'h0;
wire	[31:0]	mux_u116;
wire	[15:0]	mux_u117_u0;
wire		or_u391_u0;
reg		reg_7d7b376c_u0=1'h0;
reg		reg_7d7b376c_result_delayed_u0=1'h0;
reg	[15:0]	syncEnable_u107_u0=16'h0;
reg		reg_7d7b376c_result_delayed_result_delayed_u0=1'h0;
assign and_u1457_u0=GO&port_109251b1_;
assign and_u1458_u0=GO&port_1b0c101d_;
assign add=port_42420f9a_+32'h2;
assign and_u1459_u0=reg_712a5581_u0&port_463aad8f_;
assign or_u389_u0=and_u1459_u0|RESET;
always @(posedge CLK or posedge reg_7d7b376c_u0 or posedge or_u389_u0)
begin
if (or_u389_u0)
reg_712a5581_u0<=1'h0;
else if (reg_7d7b376c_u0)
reg_712a5581_u0<=1'h1;
else reg_712a5581_u0<=reg_712a5581_u0;
end
assign or_u390_u0=and_u1460_u0|RESET;
assign and_u1460_u0=reg_19ab1be5_u0&port_463aad8f_;
always @(posedge CLK or posedge reg_7d7b376c_result_delayed_u0 or posedge or_u390_u0)
begin
if (or_u390_u0)
reg_19ab1be5_u0<=1'h0;
else if (reg_7d7b376c_result_delayed_u0)
reg_19ab1be5_u0<=1'h1;
else reg_19ab1be5_u0<=reg_19ab1be5_u0;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u106<=port_735ece5a_;
end
assign mux_u116=(reg_7d7b376c_u0)?32'h0:32'h1;
assign mux_u117_u0=(reg_7d7b376c_u0)?syncEnable_u107_u0:syncEnable_u106;
assign or_u391_u0=reg_7d7b376c_u0|reg_7d7b376c_result_delayed_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7d7b376c_u0<=1'h0;
else reg_7d7b376c_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7d7b376c_result_delayed_u0<=1'h0;
else reg_7d7b376c_result_delayed_u0<=reg_7d7b376c_u0;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u107_u0<=port_2f0a27cf_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7d7b376c_result_delayed_result_delayed_u0<=1'h0;
else reg_7d7b376c_result_delayed_result_delayed_u0<=reg_7d7b376c_result_delayed_u0;
end
assign RESULT=GO;
assign RESULT_u862=add;
assign RESULT_u863=GO;
assign RESULT_u864=32'h1;
assign RESULT_u865=3'h1;
assign RESULT_u866=GO;
assign RESULT_u867=32'h0;
assign RESULT_u868=3'h1;
assign RESULT_u869=or_u391_u0;
assign RESULT_u870={31'b0, mux_u116[0]};
assign RESULT_u871=mux_u117_u0;
assign RESULT_u872=3'h1;
assign DONE=reg_7d7b376c_result_delayed_result_delayed_u0;
endmodule



module LL1_iunzip_stateVar_midPoint(bus_728f42fb_, bus_20ca5157_, bus_036aef22_, bus_794845ef_, bus_36d74eeb_, bus_51440103_, bus_3a6cc6f4_, bus_63d56c2a_, bus_0a115faf_, bus_110dbdeb_, bus_4867c789_);
input		bus_728f42fb_;
input		bus_20ca5157_;
input		bus_036aef22_;
input		bus_794845ef_;
input		bus_36d74eeb_;
input		bus_51440103_;
input		bus_3a6cc6f4_;
input		bus_63d56c2a_;
input		bus_0a115faf_;
input		bus_110dbdeb_;
output		bus_4867c789_;
reg		stateVar_midPoint_u1=1'h1;
wire		or_3eb4c9bf_u0;
always @(posedge bus_728f42fb_ or posedge bus_20ca5157_)
begin
if (bus_20ca5157_)
stateVar_midPoint_u1<=1'h1;
else if (or_3eb4c9bf_u0)
stateVar_midPoint_u1<=1'h0;
end
assign bus_4867c789_=stateVar_midPoint_u1;
assign or_3eb4c9bf_u0=bus_036aef22_|bus_36d74eeb_|bus_3a6cc6f4_|bus_0a115faf_;
endmodule



module LL1_iunzip_forge_memory_2x16_10(CLK, ENA, WEA, DINA, ENB, ADDRA, ADDRB, DOUTA, DOUTB, DONEA, DONEB);
input		CLK;
input		ENA;
input		WEA;
input	[15:0]	DINA;
input		ENB;
input	[31:0]	ADDRA;
input	[31:0]	ADDRB;
output	[15:0]	DOUTA;
output	[15:0]	DOUTB;
output		DONEA;
output		DONEB;
wire		wea_0;
wire	[15:0]	pre_douta_0;
wire	[15:0]	pre_doutb_0;
reg		wea_done;
reg		rea_done;
reg	[15:0]	mux_outa;
reg	[15:0]	mux_outb;
assign wea_0=WEA;
always @(posedge CLK)
begin
wea_done<=WEA;
end
assign DONEA=rea_done|wea_done;
always @(posedge CLK)
begin
end
assign DONEB=ENB;
always @(pre_douta_0)
begin
mux_outa<=pre_douta_0;
end
assign DOUTA=mux_outa;
always @(pre_doutb_0)
begin
mux_outb<=pre_doutb_0;
end
assign DOUTB=mux_outb;
// Memory array element: COL: 0, ROW: 0
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_32(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[0]), .SPO(pre_douta_0[0]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[0]));
// Memory array element: COL: 0, ROW: 1
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_33(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[1]), .SPO(pre_douta_0[1]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[1]));
// Memory array element: COL: 0, ROW: 2
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_34(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[2]), .SPO(pre_douta_0[2]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[2]));
// Memory array element: COL: 0, ROW: 3
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_35(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[3]), .SPO(pre_douta_0[3]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[3]));
// Memory array element: COL: 0, ROW: 4
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_36(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[4]), .SPO(pre_douta_0[4]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[4]));
// Memory array element: COL: 0, ROW: 5
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_37(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[5]), .SPO(pre_douta_0[5]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[5]));
// Memory array element: COL: 0, ROW: 6
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_38(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[6]), .SPO(pre_douta_0[6]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[6]));
// Memory array element: COL: 0, ROW: 7
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_39(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[7]), .SPO(pre_douta_0[7]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[7]));
// Memory array element: COL: 0, ROW: 8
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_40(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[8]), .SPO(pre_douta_0[8]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[8]));
// Memory array element: COL: 0, ROW: 9
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_41(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[9]), .SPO(pre_douta_0[9]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[9]));
// Memory array element: COL: 0, ROW: 10
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_42(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[10]), .SPO(pre_douta_0[10]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[10]));
// Memory array element: COL: 0, ROW: 11
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_43(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[11]), .SPO(pre_douta_0[11]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[11]));
// Memory array element: COL: 0, ROW: 12
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_44(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[12]), .SPO(pre_douta_0[12]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[12]));
// Memory array element: COL: 0, ROW: 13
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_45(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[13]), .SPO(pre_douta_0[13]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[13]));
// Memory array element: COL: 0, ROW: 14
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_46(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[14]), .SPO(pre_douta_0[14]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[14]));
// Memory array element: COL: 0, ROW: 15
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_47(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[15]), .SPO(pre_douta_0[15]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[15]));
endmodule



module LL1_iunzip_structuralmemory_199cf187_(CLK_u4, bus_5451230e_, bus_71688263_, bus_7304c986_, bus_3e8fafd7_, bus_4e7a128c_, bus_069ded29_, bus_016e515e_, bus_261f279e_, bus_2558522d_, bus_41de6c42_, bus_15790327_, bus_55100efa_, bus_338070be_);
input		CLK_u4;
input		bus_5451230e_;
input	[31:0]	bus_71688263_;
input	[2:0]	bus_7304c986_;
input		bus_3e8fafd7_;
input	[31:0]	bus_4e7a128c_;
input	[2:0]	bus_069ded29_;
input		bus_016e515e_;
input		bus_261f279e_;
input	[15:0]	bus_2558522d_;
output	[15:0]	bus_41de6c42_;
output		bus_15790327_;
output	[15:0]	bus_55100efa_;
output		bus_338070be_;
wire		or_2b592b1a_u0;
reg		logicalMem_8000f5b_we_delay0_u0=1'h0;
wire		not_754d82a8_u0;
wire	[15:0]	bus_5211afe3_;
wire	[15:0]	bus_23d2276f_;
wire		and_4a552b2e_u0;
wire		or_597fb922_u0;
assign or_2b592b1a_u0=bus_016e515e_|bus_261f279e_;
always @(posedge CLK_u4 or posedge bus_5451230e_)
begin
if (bus_5451230e_)
logicalMem_8000f5b_we_delay0_u0<=1'h0;
else logicalMem_8000f5b_we_delay0_u0<=bus_261f279e_;
end
assign not_754d82a8_u0=~bus_261f279e_;
LL1_iunzip_forge_memory_2x16_10 LL1_iunzip_forge_memory_2x16_10_instance0(.CLK(CLK_u4), 
  .ENA(or_2b592b1a_u0), .WEA(bus_261f279e_), .DINA(bus_2558522d_), .ADDRA(bus_4e7a128c_), 
  .DOUTA(bus_23d2276f_), .DONEA(), .ENB(bus_3e8fafd7_), .ADDRB(32'h1), .DOUTB(bus_5211afe3_), 
  .DONEB());
assign bus_41de6c42_=bus_5211afe3_;
assign bus_15790327_=bus_3e8fafd7_;
assign bus_55100efa_=bus_23d2276f_;
assign bus_338070be_=or_597fb922_u0;
assign and_4a552b2e_u0=bus_016e515e_&not_754d82a8_u0;
assign or_597fb922_u0=and_4a552b2e_u0|logicalMem_8000f5b_we_delay0_u0;
endmodule



module LL1_iunzip_streamEndFun2(CLK, RESET, GO, port_3f8bef0c_, port_3c3e7cb8_, port_74b582d8_, port_59348860_, port_38c4f7d8_, RESULT, RESULT_u873, RESULT_u874, RESULT_u875, RESULT_u876, RESULT_u877, RESULT_u878, RESULT_u879, RESULT_u880, RESULT_u881, RESULT_u882, RESULT_u883, RESULT_u884, RESULT_u885, DONE);
input		CLK;
input		RESET;
input		GO;
input		port_3f8bef0c_;
input		port_3c3e7cb8_;
input	[15:0]	port_74b582d8_;
input		port_59348860_;
input	[15:0]	port_38c4f7d8_;
output		RESULT;
output		RESULT_u873;
output		RESULT_u874;
output	[31:0]	RESULT_u875;
output	[2:0]	RESULT_u876;
output		RESULT_u877;
output	[31:0]	RESULT_u878;
output	[2:0]	RESULT_u879;
output	[15:0]	RESULT_u880;
output		RESULT_u881;
output	[15:0]	RESULT_u882;
output	[15:0]	RESULT_u883;
output	[15:0]	RESULT_u884;
output		RESULT_u885;
output		DONE;
wire	[31:0]	add;
wire		and_u1461_u0;
wire	[8:0]	subtract;
wire signed	[8:0]	greaterThanEqualTo_b_signed;
wire signed	[8:0]	greaterThanEqualTo_a_signed;
wire		greaterThanEqualTo;
wire		and_u1462_u0;
wire		not_u281_u0;
wire		and_u1463_u0;
wire	[8:0]	subtract_u8;
wire	[8:0]	mux_u118;
wire		and_u1464_u0;
wire		and_u1465_u0;
wire	[31:0]	add_u40;
wire		and_u1466_u0;
wire		and_u1468_u0;
wire	[16:0]	add_u41;
wire	[15:0]	add_u42;
wire	[15:0]	simplePinWrite;
wire		simplePinWrite_u245;
wire	[15:0]	simplePinWrite_u246;
wire	[15:0]	simplePinWrite_u247;
wire	[15:0]	simplePinWrite_u248;
wire		simplePinWrite_u249;
reg		reg_52856c80_u0=1'h0;
reg		reg_7ee62174_u0=1'h0;
reg	[31:0]	syncEnable_u108=32'h0;
wire	[31:0]	mux_u119_u0;
wire		or_u392_u0;
reg	[31:0]	syncEnable_u109_u0=32'h0;
reg	[15:0]	syncEnable_u110_u0=16'h0;
reg	[15:0]	syncEnable_u111_u0=16'h0;
assign add={31'b0, port_3f8bef0c_}+32'h0;
assign and_u1461_u0=reg_7ee62174_u0&port_3c3e7cb8_;
assign subtract={8'b0, port_3f8bef0c_}-9'h1;
assign greaterThanEqualTo_a_signed={subtract[2], subtract[2], subtract[2], subtract[2], subtract[2], subtract[2], subtract[2:0]};
assign greaterThanEqualTo_b_signed=9'h0;
assign greaterThanEqualTo=greaterThanEqualTo_a_signed>=greaterThanEqualTo_b_signed;
assign and_u1462_u0=GO&not_u281_u0;
assign not_u281_u0=~greaterThanEqualTo;
assign and_u1463_u0=GO&greaterThanEqualTo;
assign subtract_u8={8'b0, port_3f8bef0c_}-9'h1;
assign mux_u118=(and_u1465_u0)?{subtract_u8[2], subtract_u8[2], subtract_u8[2], subtract_u8[2], subtract_u8[2], subtract_u8[2], subtract_u8[2:0]}:9'h2;
assign and_u1464_u0=and_u1462_u0&GO;
assign and_u1465_u0=and_u1463_u0&GO;
assign add_u40={mux_u118[2], mux_u118[2], mux_u118[2], mux_u118[2], mux_u118[2], mux_u118[2], mux_u118[2], mux_u118[2], mux_u118[2], mux_u118[2], mux_u118[2], mux_u118[2], mux_u118[2], mux_u118[2], mux_u118[2], mux_u118[2], mux_u118[2], mux_u118[2], mux_u118[2], mux_u118[2], mux_u118[2], mux_u118[2], mux_u118[2], mux_u118[2], mux_u118[2], mux_u118[2], mux_u118[2], mux_u118[2], mux_u118[2], mux_u118[2:0]}+32'h0;
assign and_u1466_u0=reg_7ee62174_u0&port_59348860_;
assign and_u1468_u0=reg_52856c80_u0&port_3c3e7cb8_;
assign add_u41={syncEnable_u111_u0[15], syncEnable_u111_u0}+{port_74b582d8_[15], port_74b582d8_};
assign add_u42=syncEnable_u110_u0+{add_u41[16], add_u41[16:2]};
assign simplePinWrite=add_u42&{16{reg_52856c80_u0}};
assign simplePinWrite_u245=reg_52856c80_u0&{1{reg_52856c80_u0}};
assign simplePinWrite_u246=16'h1&{16{1'h1}};
assign simplePinWrite_u247=16'h1&{16{1'h1}};
assign simplePinWrite_u248=add_u42&{16{reg_52856c80_u0}};
assign simplePinWrite_u249=reg_52856c80_u0&{1{reg_52856c80_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_52856c80_u0<=1'h0;
else reg_52856c80_u0<=reg_7ee62174_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7ee62174_u0<=1'h0;
else reg_7ee62174_u0<=GO;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u108<={add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2:0]};
end
assign mux_u119_u0=(reg_7ee62174_u0)?syncEnable_u108:32'h0;
assign or_u392_u0=reg_7ee62174_u0|reg_52856c80_u0;
always @(posedge CLK)
begin
if (GO)
syncEnable_u109_u0<=add_u40;
end
always @(posedge CLK)
begin
if (reg_7ee62174_u0)
syncEnable_u110_u0<=port_74b582d8_;
end
always @(posedge CLK)
begin
if (reg_7ee62174_u0)
syncEnable_u111_u0<=port_38c4f7d8_;
end
assign RESULT=GO;
assign RESULT_u873=1'h0;
assign RESULT_u874=or_u392_u0;
assign RESULT_u875=mux_u119_u0;
assign RESULT_u876=3'h1;
assign RESULT_u877=reg_7ee62174_u0;
assign RESULT_u878=syncEnable_u109_u0;
assign RESULT_u879=3'h1;
assign RESULT_u880=simplePinWrite_u248;
assign RESULT_u881=simplePinWrite_u245;
assign RESULT_u882=simplePinWrite;
assign RESULT_u883=simplePinWrite_u246;
assign RESULT_u884=simplePinWrite_u247;
assign RESULT_u885=simplePinWrite_u249;
assign DONE=reg_52856c80_u0;
endmodule



module LL1_iunzip_Kicker_26(CLK, RESET, bus_251f35c9_);
input		CLK;
input		RESET;
output		bus_251f35c9_;
wire		bus_7d86fec0_;
wire		bus_3e801401_;
wire		bus_19c5edac_;
reg		kicker_2=1'h0;
reg		kicker_1=1'h0;
reg		kicker_res=1'h0;
wire		bus_68ea3357_;
assign bus_7d86fec0_=bus_19c5edac_&kicker_1;
assign bus_3e801401_=kicker_1&bus_19c5edac_&bus_68ea3357_;
assign bus_19c5edac_=~RESET;
always @(posedge CLK)
begin
kicker_2<=bus_7d86fec0_;
end
always @(posedge CLK)
begin
kicker_1<=bus_19c5edac_;
end
assign bus_251f35c9_=kicker_res;
always @(posedge CLK)
begin
kicker_res<=bus_3e801401_;
end
assign bus_68ea3357_=~kicker_2;
endmodule



module LL1_iunzip_simplememoryreferee_52a82a09_(bus_2453e19e_, bus_1b3c311c_, bus_06bb3bca_, bus_7f823762_, bus_33f699d7_, bus_0e87d9ae_, bus_51e962ad_, bus_43cb9bbb_, bus_5be4b948_, bus_238bf419_, bus_7bd172a7_, bus_0319de32_, bus_60a35d69_, bus_7475072e_, bus_7cd5d094_, bus_2e6c9d65_, bus_735b4165_, bus_2da416ce_, bus_455d1534_, bus_5347953e_, bus_1ebd7ee4_, bus_707f0c59_, bus_1ec36984_, bus_5239f197_, bus_11305c14_, bus_2a9ec1c5_, bus_578aeeb2_, bus_17d4c247_, bus_1d3e0f48_, bus_26f430ba_, bus_5c92336e_, bus_69d30eb5_, bus_05a209b3_, bus_4f3b4ae4_, bus_50a40b11_, bus_167013f4_, bus_66064e11_, bus_71da01b9_);
input		bus_2453e19e_;
input		bus_1b3c311c_;
input		bus_06bb3bca_;
input	[15:0]	bus_7f823762_;
input		bus_33f699d7_;
input	[15:0]	bus_0e87d9ae_;
input	[31:0]	bus_51e962ad_;
input	[2:0]	bus_43cb9bbb_;
input		bus_5be4b948_;
input		bus_238bf419_;
input	[15:0]	bus_7bd172a7_;
input	[31:0]	bus_0319de32_;
input	[2:0]	bus_60a35d69_;
input		bus_7475072e_;
input		bus_7cd5d094_;
input	[15:0]	bus_2e6c9d65_;
input	[31:0]	bus_735b4165_;
input	[2:0]	bus_2da416ce_;
input		bus_455d1534_;
input	[31:0]	bus_5347953e_;
input	[2:0]	bus_1ebd7ee4_;
input		bus_707f0c59_;
input	[31:0]	bus_1ec36984_;
input	[2:0]	bus_5239f197_;
output	[15:0]	bus_11305c14_;
output	[31:0]	bus_2a9ec1c5_;
output		bus_578aeeb2_;
output		bus_17d4c247_;
output	[2:0]	bus_1d3e0f48_;
output		bus_26f430ba_;
output	[15:0]	bus_5c92336e_;
output		bus_69d30eb5_;
output	[15:0]	bus_05a209b3_;
output		bus_4f3b4ae4_;
output	[15:0]	bus_50a40b11_;
output		bus_167013f4_;
output	[15:0]	bus_66064e11_;
output		bus_71da01b9_;
reg		done_qual_u55_u0=1'h0;
wire		not_66f52031_u0;
wire		not_15d5b152_u0;
wire	[31:0]	mux_01442848_u0;
reg		done_qual_u56_u0=1'h0;
wire		or_3d932703_u0;
wire		and_70be256e_u0;
wire		or_18a2cdb3_u0;
wire		not_187827e9_u0;
wire		and_17fe43a9_u0;
wire		not_20d9cbce_u0;
wire		not_035f2b45_u0;
wire		and_6b4acc50_u0;
wire		or_7bf24c2e_u0;
wire		or_694641db_u0;
wire		or_6cc5e89b_u0;
wire		or_33c2389c_u0;
wire		and_7ea02ffe_u0;
reg		done_qual_u57_u0=1'h0;
wire	[15:0]	mux_302170cc_u0;
wire		or_5151513c_u0;
wire		or_4a02aaac_u0;
reg		done_qual_u58_u0=1'h0;
wire		and_57de3d6f_u0;
reg		done_qual_u59_u0=1'h0;
wire		or_260eab74_u0;
always @(posedge bus_2453e19e_)
begin
if (bus_1b3c311c_)
done_qual_u55_u0<=1'h0;
else done_qual_u55_u0<=or_18a2cdb3_u0;
end
assign not_66f52031_u0=~bus_06bb3bca_;
assign not_15d5b152_u0=~bus_06bb3bca_;
assign mux_01442848_u0=({32{bus_33f699d7_}}&{31'b0, bus_51e962ad_[0]})|({32{or_18a2cdb3_u0}}&bus_0319de32_)|({32{or_694641db_u0}}&bus_735b4165_)|({32{bus_455d1534_}}&bus_5347953e_)|({32{bus_707f0c59_}}&bus_1ec36984_);
always @(posedge bus_2453e19e_)
begin
if (bus_1b3c311c_)
done_qual_u56_u0<=1'h0;
else done_qual_u56_u0<=bus_455d1534_;
end
assign or_3d932703_u0=bus_33f699d7_|done_qual_u57_u0;
assign and_70be256e_u0=or_33c2389c_u0&bus_06bb3bca_;
assign or_18a2cdb3_u0=bus_5be4b948_|bus_238bf419_;
assign not_187827e9_u0=~bus_06bb3bca_;
assign and_17fe43a9_u0=or_3d932703_u0&bus_06bb3bca_;
assign not_20d9cbce_u0=~bus_06bb3bca_;
assign not_035f2b45_u0=~bus_06bb3bca_;
assign and_6b4acc50_u0=or_5151513c_u0&bus_06bb3bca_;
assign or_7bf24c2e_u0=bus_707f0c59_|done_qual_u59_u0;
assign or_694641db_u0=bus_7475072e_|bus_7cd5d094_;
assign or_6cc5e89b_u0=or_18a2cdb3_u0|done_qual_u55_u0;
assign or_33c2389c_u0=bus_455d1534_|done_qual_u56_u0;
assign and_7ea02ffe_u0=or_7bf24c2e_u0&bus_06bb3bca_;
always @(posedge bus_2453e19e_)
begin
if (bus_1b3c311c_)
done_qual_u57_u0<=1'h0;
else done_qual_u57_u0<=bus_33f699d7_;
end
assign mux_302170cc_u0=({16{bus_33f699d7_}}&bus_0e87d9ae_)|({16{bus_238bf419_}}&bus_7bd172a7_)|({16{bus_7cd5d094_}}&bus_2e6c9d65_);
assign or_5151513c_u0=or_694641db_u0|done_qual_u58_u0;
assign or_4a02aaac_u0=bus_33f699d7_|bus_238bf419_|bus_7cd5d094_;
always @(posedge bus_2453e19e_)
begin
if (bus_1b3c311c_)
done_qual_u58_u0<=1'h0;
else done_qual_u58_u0<=or_694641db_u0;
end
assign bus_11305c14_=mux_302170cc_u0;
assign bus_2a9ec1c5_=mux_01442848_u0;
assign bus_578aeeb2_=or_4a02aaac_u0;
assign bus_17d4c247_=or_260eab74_u0;
assign bus_1d3e0f48_=3'h1;
assign bus_26f430ba_=and_17fe43a9_u0;
assign bus_5c92336e_=bus_7f823762_;
assign bus_69d30eb5_=and_57de3d6f_u0;
assign bus_05a209b3_=bus_7f823762_;
assign bus_4f3b4ae4_=and_6b4acc50_u0;
assign bus_50a40b11_=bus_7f823762_;
assign bus_167013f4_=and_70be256e_u0;
assign bus_66064e11_=bus_7f823762_;
assign bus_71da01b9_=and_7ea02ffe_u0;
assign and_57de3d6f_u0=or_6cc5e89b_u0&bus_06bb3bca_;
always @(posedge bus_2453e19e_)
begin
if (bus_1b3c311c_)
done_qual_u59_u0<=1'h0;
else done_qual_u59_u0<=bus_707f0c59_;
end
assign or_260eab74_u0=bus_33f699d7_|or_18a2cdb3_u0|or_694641db_u0|bus_455d1534_|bus_707f0c59_;
endmodule



module LL1_iunzip_streamFun2(CLK, RESET, GO, port_4b4b2561_, port_5a2a759b_, port_741f83f2_, port_3d5a0933_, port_6091a1b3_, port_3f9a965b_, port_15d252f1_, port_189d0bed_, RESULT, RESULT_u886, RESULT_u887, RESULT_u888, RESULT_u889, RESULT_u890, RESULT_u891, RESULT_u892, RESULT_u893, RESULT_u894, RESULT_u895, RESULT_u896, RESULT_u897, RESULT_u898, RESULT_u899, RESULT_u900, RESULT_u901, RESULT_u902, DONE);
input		CLK;
input		RESET;
input		GO;
input		port_4b4b2561_;
input	[31:0]	port_5a2a759b_;
input		port_741f83f2_;
input	[15:0]	port_3d5a0933_;
input		port_6091a1b3_;
input	[15:0]	port_3f9a965b_;
input		port_15d252f1_;
input	[15:0]	port_189d0bed_;
output		RESULT;
output		RESULT_u886;
output		RESULT_u887;
output	[31:0]	RESULT_u888;
output		RESULT_u889;
output	[31:0]	RESULT_u890;
output	[2:0]	RESULT_u891;
output		RESULT_u892;
output	[31:0]	RESULT_u893;
output	[2:0]	RESULT_u894;
output		RESULT_u895;
output	[31:0]	RESULT_u896;
output	[15:0]	RESULT_u897;
output	[2:0]	RESULT_u898;
output		RESULT_u899;
output	[15:0]	RESULT_u900;
output	[15:0]	RESULT_u901;
output		RESULT_u902;
output		DONE;
wire		simplePinWrite;
reg		reg_33b75493_u0=1'h0;
wire		and_u1471_u0;
wire		or_u393_u0;
wire	[31:0]	add;
wire		and_u1472_u0;
wire	[8:0]	subtract;
wire signed	[8:0]	greaterThanEqualTo_a_signed;
wire signed	[8:0]	greaterThanEqualTo_b_signed;
wire		greaterThanEqualTo;
wire		and_u1473_u0;
wire		not_u282_u0;
wire		and_u1474_u0;
wire	[8:0]	subtract_u9;
wire	[8:0]	mux_u120;
wire		and_u1475_u0;
wire		and_u1476_u0;
wire	[31:0]	add_u43;
wire		and_u1477_u0;
wire		and_u1479_u0;
wire	[16:0]	add_u44;
wire	[15:0]	add_u45;
wire	[31:0]	add_u46;
wire	[15:0]	simplePinWrite_u250;
wire	[15:0]	simplePinWrite_u251;
wire		simplePinWrite_u252;
reg		reg_4c8cff89_u0=1'h0;
wire	[31:0]	mux_u121_u0;
wire		or_u394_u0;
wire	[31:0]	mux_u122_u0;
reg	[31:0]	syncEnable_u112=32'h0;
reg	[15:0]	syncEnable_u113_u0=16'h0;
reg	[31:0]	syncEnable_u114_u0=32'h0;
reg		reg_4c8cff89_result_delayed_u0=1'h0;
reg		reg_43c7d006_u0=1'h0;
reg	[15:0]	syncEnable_u115_u0=16'h0;
reg	[15:0]	syncEnable_u116_u0=16'h0;
assign simplePinWrite=GO&{1{GO}};
always @(posedge CLK or posedge reg_43c7d006_u0 or posedge or_u393_u0)
begin
if (or_u393_u0)
reg_33b75493_u0<=1'h0;
else if (reg_43c7d006_u0)
reg_33b75493_u0<=1'h1;
else reg_33b75493_u0<=reg_33b75493_u0;
end
assign and_u1471_u0=reg_33b75493_u0&port_15d252f1_;
assign or_u393_u0=and_u1471_u0|RESET;
assign add={31'b0, port_4b4b2561_}+32'h0;
assign and_u1472_u0=reg_4c8cff89_u0&port_741f83f2_;
assign subtract={8'b0, port_4b4b2561_}-9'h1;
assign greaterThanEqualTo_a_signed={subtract[2], subtract[2], subtract[2], subtract[2], subtract[2], subtract[2], subtract[2:0]};
assign greaterThanEqualTo_b_signed=9'h0;
assign greaterThanEqualTo=greaterThanEqualTo_a_signed>=greaterThanEqualTo_b_signed;
assign and_u1473_u0=GO&not_u282_u0;
assign not_u282_u0=~greaterThanEqualTo;
assign and_u1474_u0=GO&greaterThanEqualTo;
assign subtract_u9={8'b0, port_4b4b2561_}-9'h1;
assign mux_u120=(and_u1476_u0)?{subtract_u9[2], subtract_u9[2], subtract_u9[2], subtract_u9[2], subtract_u9[2], subtract_u9[2], subtract_u9[2:0]}:9'h2;
assign and_u1475_u0=and_u1473_u0&GO;
assign and_u1476_u0=and_u1474_u0&GO;
assign add_u43={mux_u120[2], mux_u120[2], mux_u120[2], mux_u120[2], mux_u120[2], mux_u120[2], mux_u120[2], mux_u120[2], mux_u120[2], mux_u120[2], mux_u120[2], mux_u120[2], mux_u120[2], mux_u120[2], mux_u120[2], mux_u120[2], mux_u120[2], mux_u120[2], mux_u120[2], mux_u120[2], mux_u120[2], mux_u120[2], mux_u120[2], mux_u120[2], mux_u120[2], mux_u120[2], mux_u120[2], mux_u120[2], mux_u120[2], mux_u120[2:0]}+32'h0;
assign and_u1477_u0=reg_4c8cff89_u0&port_15d252f1_;
assign and_u1479_u0=reg_4c8cff89_result_delayed_u0&port_741f83f2_;
assign add_u44={syncEnable_u116_u0[15], syncEnable_u116_u0}+{port_3d5a0933_[15], port_3d5a0933_};
assign add_u45=syncEnable_u113_u0+{add_u44[16], add_u44[16:2]};
assign add_u46=port_5a2a759b_+32'h1;
assign simplePinWrite_u250=add_u45&{16{reg_4c8cff89_result_delayed_u0}};
assign simplePinWrite_u251=16'h1&{16{1'h1}};
assign simplePinWrite_u252=reg_4c8cff89_result_delayed_u0&{1{reg_4c8cff89_result_delayed_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4c8cff89_u0<=1'h0;
else reg_4c8cff89_u0<=reg_43c7d006_u0;
end
assign mux_u121_u0=(reg_43c7d006_u0)?32'h0:syncEnable_u112;
assign or_u394_u0=reg_4c8cff89_u0|reg_4c8cff89_result_delayed_u0;
assign mux_u122_u0=(reg_4c8cff89_u0)?syncEnable_u114_u0:32'h0;
always @(posedge CLK)
begin
if (GO)
syncEnable_u112<=add_u43;
end
always @(posedge CLK)
begin
if (reg_4c8cff89_u0)
syncEnable_u113_u0<=port_3d5a0933_;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u114_u0<={add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2:0]};
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4c8cff89_result_delayed_u0<=1'h0;
else reg_4c8cff89_result_delayed_u0<=reg_4c8cff89_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_43c7d006_u0<=1'h0;
else reg_43c7d006_u0<=GO;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u115_u0<=port_189d0bed_;
end
always @(posedge CLK)
begin
if (reg_4c8cff89_u0)
syncEnable_u116_u0<=port_3f9a965b_;
end
assign RESULT=GO;
assign RESULT_u886=1'h0;
assign RESULT_u887=GO;
assign RESULT_u888=add_u46;
assign RESULT_u889=or_u394_u0;
assign RESULT_u890=mux_u122_u0;
assign RESULT_u891=3'h1;
assign RESULT_u892=reg_4c8cff89_u0;
assign RESULT_u893=mux_u121_u0;
assign RESULT_u894=3'h1;
assign RESULT_u895=reg_43c7d006_u0;
assign RESULT_u896=mux_u121_u0;
assign RESULT_u897=syncEnable_u115_u0;
assign RESULT_u898=3'h1;
assign RESULT_u899=simplePinWrite;
assign RESULT_u900=simplePinWrite_u250;
assign RESULT_u901=simplePinWrite_u251;
assign RESULT_u902=simplePinWrite_u252;
assign DONE=reg_4c8cff89_result_delayed_u0;
endmodule



module LL1_iunzip_endianswapper_3216ffed_(endianswapper_3216ffed_in, endianswapper_3216ffed_out);
input	[1:0]	endianswapper_3216ffed_in;
output	[1:0]	endianswapper_3216ffed_out;
assign endianswapper_3216ffed_out=endianswapper_3216ffed_in;
endmodule



module LL1_iunzip_endianswapper_258e9931_(endianswapper_258e9931_in, endianswapper_258e9931_out);
input	[1:0]	endianswapper_258e9931_in;
output	[1:0]	endianswapper_258e9931_out;
assign endianswapper_258e9931_out=endianswapper_258e9931_in;
endmodule



module LL1_iunzip_stateVar_fsmOldState_LL1_iunzip(bus_20ec10f4_, bus_09f76d0f_, bus_7508f03a_, bus_078eb971_, bus_7d60e04a_);
input		bus_20ec10f4_;
input		bus_09f76d0f_;
input		bus_7508f03a_;
input	[1:0]	bus_078eb971_;
output	[1:0]	bus_7d60e04a_;
reg	[1:0]	stateVar_fsmOldState_LL1_iunzip_u0=2'h0;
wire	[1:0]	endianswapper_3216ffed_out;
wire	[1:0]	endianswapper_258e9931_out;
always @(posedge bus_20ec10f4_ or posedge bus_09f76d0f_)
begin
if (bus_09f76d0f_)
stateVar_fsmOldState_LL1_iunzip_u0<=2'h0;
else if (bus_7508f03a_)
stateVar_fsmOldState_LL1_iunzip_u0<=endianswapper_3216ffed_out;
end
assign bus_7d60e04a_=endianswapper_258e9931_out;
LL1_iunzip_endianswapper_3216ffed_ LL1_iunzip_endianswapper_3216ffed__1(.endianswapper_3216ffed_in(bus_078eb971_), 
  .endianswapper_3216ffed_out(endianswapper_3216ffed_out));
LL1_iunzip_endianswapper_258e9931_ LL1_iunzip_endianswapper_258e9931__1(.endianswapper_258e9931_in(stateVar_fsmOldState_LL1_iunzip_u0), 
  .endianswapper_258e9931_out(endianswapper_258e9931_out));
endmodule



module LL1_iunzip_simplememoryreferee_7e53def4_(bus_5e9a9b98_, bus_0b4a27a7_, bus_6ceb0c3b_, bus_3ec3c7a3_, bus_50a4ddaf_, bus_04a67922_, bus_40e70fc3_, bus_5a00092e_, bus_38e2b04c_, bus_422fb56c_, bus_732498ad_, bus_306ebd50_, bus_15657ed6_, bus_7e9b0677_);
input		bus_5e9a9b98_;
input		bus_0b4a27a7_;
input		bus_6ceb0c3b_;
input	[15:0]	bus_3ec3c7a3_;
input		bus_50a4ddaf_;
input	[31:0]	bus_04a67922_;
input	[2:0]	bus_40e70fc3_;
output	[15:0]	bus_5a00092e_;
output	[31:0]	bus_38e2b04c_;
output		bus_422fb56c_;
output		bus_732498ad_;
output	[2:0]	bus_306ebd50_;
output	[15:0]	bus_15657ed6_;
output		bus_7e9b0677_;
assign bus_5a00092e_=16'h0;
assign bus_38e2b04c_=32'h1;
assign bus_422fb56c_=1'h0;
assign bus_732498ad_=bus_50a4ddaf_;
assign bus_306ebd50_=3'h1;
assign bus_15657ed6_=bus_3ec3c7a3_;
assign bus_7e9b0677_=bus_6ceb0c3b_;
endmodule



module LL1_iunzip_stateVar_In1PortEnable(bus_482b48c2_, bus_414ca731_, bus_27b57e02_, bus_119b13c9_, bus_26b0e73f_);
input		bus_482b48c2_;
input		bus_414ca731_;
input		bus_27b57e02_;
input		bus_119b13c9_;
output		bus_26b0e73f_;
reg		stateVar_In1PortEnable_u1=1'h0;
assign bus_26b0e73f_=stateVar_In1PortEnable_u1;
always @(posedge bus_482b48c2_ or posedge bus_414ca731_)
begin
if (bus_414ca731_)
stateVar_In1PortEnable_u1<=1'h0;
else if (bus_27b57e02_)
stateVar_In1PortEnable_u1<=bus_119b13c9_;
end
endmodule



module LL1_iunzip_endianswapper_101754b7_(endianswapper_101754b7_in, endianswapper_101754b7_out);
input	[1:0]	endianswapper_101754b7_in;
output	[1:0]	endianswapper_101754b7_out;
assign endianswapper_101754b7_out=endianswapper_101754b7_in;
endmodule



module LL1_iunzip_endianswapper_0b341926_(endianswapper_0b341926_in, endianswapper_0b341926_out);
input	[1:0]	endianswapper_0b341926_in;
output	[1:0]	endianswapper_0b341926_out;
assign endianswapper_0b341926_out=endianswapper_0b341926_in;
endmodule



module LL1_iunzip_stateVar_fsmState_LL1_iunzip(bus_781a7383_, bus_11069aeb_, bus_2457321f_, bus_2a0ed9bb_, bus_3c6b3bea_);
input		bus_781a7383_;
input		bus_11069aeb_;
input		bus_2457321f_;
input	[1:0]	bus_2a0ed9bb_;
output	[1:0]	bus_3c6b3bea_;
wire	[1:0]	endianswapper_101754b7_out;
wire	[1:0]	endianswapper_0b341926_out;
reg	[1:0]	stateVar_fsmState_LL1_iunzip_u0=2'h0;
LL1_iunzip_endianswapper_101754b7_ LL1_iunzip_endianswapper_101754b7__1(.endianswapper_101754b7_in(bus_2a0ed9bb_), 
  .endianswapper_101754b7_out(endianswapper_101754b7_out));
LL1_iunzip_endianswapper_0b341926_ LL1_iunzip_endianswapper_0b341926__1(.endianswapper_0b341926_in(stateVar_fsmState_LL1_iunzip_u0), 
  .endianswapper_0b341926_out(endianswapper_0b341926_out));
assign bus_3c6b3bea_=endianswapper_0b341926_out;
always @(posedge bus_781a7383_ or posedge bus_11069aeb_)
begin
if (bus_11069aeb_)
stateVar_fsmState_LL1_iunzip_u0<=2'h0;
else if (bus_2457321f_)
stateVar_fsmState_LL1_iunzip_u0<=endianswapper_101754b7_out;
end
endmodule



module LL1_iunzip_forge_memory_3x16_11(CLK, ENA, WEA, DINA, ENB, ADDRA, ADDRB, DOUTA, DOUTB, DONEA, DONEB);
input		CLK;
input		ENA;
input		WEA;
input	[15:0]	DINA;
input		ENB;
input	[31:0]	ADDRA;
input	[31:0]	ADDRB;
output	[15:0]	DOUTA;
output	[15:0]	DOUTB;
output		DONEA;
output		DONEB;
wire		wea_0;
wire	[15:0]	pre_douta_0;
wire	[15:0]	pre_doutb_0;
reg		wea_done;
reg		rea_done;
reg	[15:0]	mux_outa;
reg	[15:0]	mux_outb;
assign wea_0=WEA;
always @(posedge CLK)
begin
wea_done<=WEA;
end
assign DONEA=rea_done|wea_done;
always @(posedge CLK)
begin
end
assign DONEB=ENB;
always @(pre_douta_0)
begin
mux_outa<=pre_douta_0;
end
assign DOUTA=mux_outa;
always @(pre_doutb_0)
begin
mux_outb<=pre_doutb_0;
end
assign DOUTB=mux_outb;
// Memory array element: COL: 0, ROW: 0
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_48(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[0]), .SPO(pre_douta_0[0]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[0]));
// Memory array element: COL: 0, ROW: 1
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_49(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[1]), .SPO(pre_douta_0[1]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[1]));
// Memory array element: COL: 0, ROW: 2
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_50(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[2]), .SPO(pre_douta_0[2]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[2]));
// Memory array element: COL: 0, ROW: 3
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_51(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[3]), .SPO(pre_douta_0[3]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[3]));
// Memory array element: COL: 0, ROW: 4
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_52(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[4]), .SPO(pre_douta_0[4]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[4]));
// Memory array element: COL: 0, ROW: 5
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_53(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[5]), .SPO(pre_douta_0[5]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[5]));
// Memory array element: COL: 0, ROW: 6
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_54(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[6]), .SPO(pre_douta_0[6]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[6]));
// Memory array element: COL: 0, ROW: 7
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_55(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[7]), .SPO(pre_douta_0[7]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[7]));
// Memory array element: COL: 0, ROW: 8
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_56(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[8]), .SPO(pre_douta_0[8]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[8]));
// Memory array element: COL: 0, ROW: 9
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_57(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[9]), .SPO(pre_douta_0[9]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[9]));
// Memory array element: COL: 0, ROW: 10
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_58(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[10]), .SPO(pre_douta_0[10]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[10]));
// Memory array element: COL: 0, ROW: 11
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_59(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[11]), .SPO(pre_douta_0[11]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[11]));
// Memory array element: COL: 0, ROW: 12
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_60(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[12]), .SPO(pre_douta_0[12]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[12]));
// Memory array element: COL: 0, ROW: 13
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_61(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[13]), .SPO(pre_douta_0[13]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[13]));
// Memory array element: COL: 0, ROW: 14
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_62(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[14]), .SPO(pre_douta_0[14]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[14]));
// Memory array element: COL: 0, ROW: 15
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_63(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[15]), .SPO(pre_douta_0[15]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[15]));
endmodule



module LL1_iunzip_structuralmemory_65c92979_(CLK_u5, bus_1dee1645_, bus_36216417_, bus_06d309bc_, bus_6296f247_, bus_083d81f6_, bus_3786b3c5_, bus_0f87e737_, bus_7a6a921b_, bus_2c10caec_, bus_1deedea6_, bus_0de9df36_, bus_2c07dd11_, bus_454c7853_);
input		CLK_u5;
input		bus_1dee1645_;
input	[31:0]	bus_36216417_;
input	[2:0]	bus_06d309bc_;
input		bus_6296f247_;
input	[31:0]	bus_083d81f6_;
input	[2:0]	bus_3786b3c5_;
input		bus_0f87e737_;
input		bus_7a6a921b_;
input	[15:0]	bus_2c10caec_;
output	[15:0]	bus_1deedea6_;
output		bus_0de9df36_;
output	[15:0]	bus_2c07dd11_;
output		bus_454c7853_;
wire		not_734df1ec_u0;
wire	[15:0]	bus_6aadd3b9_;
wire	[15:0]	bus_2ac66d9e_;
wire		or_4642dc48_u0;
reg		logicalMem_31bb9af_we_delay0_u0=1'h0;
wire		and_301160c6_u0;
wire		or_4c4c6133_u0;
assign not_734df1ec_u0=~bus_7a6a921b_;
LL1_iunzip_forge_memory_3x16_11 LL1_iunzip_forge_memory_3x16_11_instance0(.CLK(CLK_u5), 
  .ENA(or_4642dc48_u0), .WEA(bus_7a6a921b_), .DINA(bus_2c10caec_), .ADDRA(bus_083d81f6_), 
  .DOUTA(bus_6aadd3b9_), .DONEA(), .ENB(bus_6296f247_), .ADDRB(bus_36216417_), .DOUTB(bus_2ac66d9e_), 
  .DONEB());
assign or_4642dc48_u0=bus_0f87e737_|bus_7a6a921b_;
always @(posedge CLK_u5 or posedge bus_1dee1645_)
begin
if (bus_1dee1645_)
logicalMem_31bb9af_we_delay0_u0<=1'h0;
else logicalMem_31bb9af_we_delay0_u0<=bus_7a6a921b_;
end
assign bus_1deedea6_=bus_2ac66d9e_;
assign bus_0de9df36_=bus_6296f247_;
assign bus_2c07dd11_=bus_6aadd3b9_;
assign bus_454c7853_=or_4c4c6133_u0;
assign and_301160c6_u0=bus_0f87e737_&not_734df1ec_u0;
assign or_4c4c6133_u0=and_301160c6_u0|logicalMem_31bb9af_we_delay0_u0;
endmodule



module LL1_iunzip_endianswapper_40d3b487_(endianswapper_40d3b487_in, endianswapper_40d3b487_out);
input	[31:0]	endianswapper_40d3b487_in;
output	[31:0]	endianswapper_40d3b487_out;
assign endianswapper_40d3b487_out=endianswapper_40d3b487_in;
endmodule



module LL1_iunzip_endianswapper_12c8575f_(endianswapper_12c8575f_in, endianswapper_12c8575f_out);
input	[31:0]	endianswapper_12c8575f_in;
output	[31:0]	endianswapper_12c8575f_out;
assign endianswapper_12c8575f_out=endianswapper_12c8575f_in;
endmodule



module LL1_iunzip_stateVar_In1TokenIndex(bus_028bcee6_, bus_3ce31b6e_, bus_3da9e3d5_, bus_4515a94c_, bus_22baa6c8_);
input		bus_028bcee6_;
input		bus_3ce31b6e_;
input		bus_3da9e3d5_;
input	[31:0]	bus_4515a94c_;
output	[31:0]	bus_22baa6c8_;
wire	[31:0]	endianswapper_40d3b487_out;
wire	[31:0]	endianswapper_12c8575f_out;
reg	[31:0]	stateVar_In1TokenIndex_u1=32'h0;
LL1_iunzip_endianswapper_40d3b487_ LL1_iunzip_endianswapper_40d3b487__1(.endianswapper_40d3b487_in(stateVar_In1TokenIndex_u1), 
  .endianswapper_40d3b487_out(endianswapper_40d3b487_out));
assign bus_22baa6c8_=endianswapper_40d3b487_out;
LL1_iunzip_endianswapper_12c8575f_ LL1_iunzip_endianswapper_12c8575f__1(.endianswapper_12c8575f_in(bus_4515a94c_), 
  .endianswapper_12c8575f_out(endianswapper_12c8575f_out));
always @(posedge bus_028bcee6_ or posedge bus_3ce31b6e_)
begin
if (bus_3ce31b6e_)
stateVar_In1TokenIndex_u1<=32'h0;
else if (bus_3da9e3d5_)
stateVar_In1TokenIndex_u1<=endianswapper_12c8575f_out;
end
endmodule



module LL1_iunzip_endianswapper_331ca0aa_(endianswapper_331ca0aa_in, endianswapper_331ca0aa_out);
input	[31:0]	endianswapper_331ca0aa_in;
output	[31:0]	endianswapper_331ca0aa_out;
assign endianswapper_331ca0aa_out=endianswapper_331ca0aa_in;
endmodule



module LL1_iunzip_endianswapper_2fd0da88_(endianswapper_2fd0da88_in, endianswapper_2fd0da88_out);
input	[31:0]	endianswapper_2fd0da88_in;
output	[31:0]	endianswapper_2fd0da88_out;
assign endianswapper_2fd0da88_out={endianswapper_2fd0da88_in[31:2], 1'b1, endianswapper_2fd0da88_in[0]};
endmodule



module LL1_iunzip_stateVar_In1MaxTokenIndex(bus_21b70cb9_, bus_0a95df40_, bus_68994182_, bus_5519f449_, bus_072b555f_);
input		bus_21b70cb9_;
input		bus_0a95df40_;
input		bus_68994182_;
input	[31:0]	bus_5519f449_;
output	[31:0]	bus_072b555f_;
wire	[31:0]	endianswapper_331ca0aa_out;
wire	[31:0]	endianswapper_2fd0da88_out;
reg	[31:0]	stateVar_In1MaxTokenIndex_u1=32'h0;
LL1_iunzip_endianswapper_331ca0aa_ LL1_iunzip_endianswapper_331ca0aa__1(.endianswapper_331ca0aa_in(stateVar_In1MaxTokenIndex_u1), 
  .endianswapper_331ca0aa_out(endianswapper_331ca0aa_out));
LL1_iunzip_endianswapper_2fd0da88_ LL1_iunzip_endianswapper_2fd0da88__1(.endianswapper_2fd0da88_in({bus_5519f449_[31:2], 1'b0, bus_5519f449_[0]}), 
  .endianswapper_2fd0da88_out(endianswapper_2fd0da88_out));
assign bus_072b555f_=endianswapper_331ca0aa_out;
always @(posedge bus_21b70cb9_ or posedge bus_0a95df40_)
begin
if (bus_0a95df40_)
stateVar_In1MaxTokenIndex_u1<=32'h0;
else if (bus_68994182_)
stateVar_In1MaxTokenIndex_u1<={endianswapper_2fd0da88_out[31:2], 1'b1, endianswapper_2fd0da88_out[0]};
end
endmodule



module LL1_iunzip_streamEndFun1(CLK, RESET, GO, port_3b9b03c5_, port_53886836_, port_63c1f3c3_, port_2d39d825_, port_768c8415_, RESULT, RESULT_u903, RESULT_u904, RESULT_u905, RESULT_u906, RESULT_u907, RESULT_u908, RESULT_u909, RESULT_u910, RESULT_u911, RESULT_u912, RESULT_u913, RESULT_u914, RESULT_u915, DONE);
input		CLK;
input		RESET;
input		GO;
input		port_3b9b03c5_;
input		port_53886836_;
input	[15:0]	port_63c1f3c3_;
input		port_2d39d825_;
input	[15:0]	port_768c8415_;
output		RESULT;
output		RESULT_u903;
output		RESULT_u904;
output	[31:0]	RESULT_u905;
output	[2:0]	RESULT_u906;
output		RESULT_u907;
output	[31:0]	RESULT_u908;
output	[2:0]	RESULT_u909;
output	[15:0]	RESULT_u910;
output		RESULT_u911;
output	[15:0]	RESULT_u912;
output	[15:0]	RESULT_u913;
output	[15:0]	RESULT_u914;
output		RESULT_u915;
output		DONE;
wire	[31:0]	add;
wire		and_u1481_u0;
wire	[8:0]	subtract;
wire signed	[8:0]	greaterThanEqualTo_b_signed;
wire signed	[8:0]	greaterThanEqualTo_a_signed;
wire		greaterThanEqualTo;
wire		and_u1482_u0;
wire		and_u1483_u0;
wire		not_u283_u0;
wire	[8:0]	subtract_u10;
wire		and_u1484_u0;
wire		and_u1485_u0;
wire	[8:0]	mux_u123;
wire	[31:0]	add_u47;
wire		and_u1486_u0;
wire		and_u1488_u0;
wire	[16:0]	add_u48;
wire	[15:0]	subtract_u11;
wire	[15:0]	simplePinWrite;
wire		simplePinWrite_u253;
wire	[15:0]	simplePinWrite_u254;
wire	[15:0]	simplePinWrite_u255;
wire		simplePinWrite_u256;
wire	[15:0]	simplePinWrite_u257;
reg	[31:0]	syncEnable_u117=32'h0;
reg	[31:0]	syncEnable_u118_u0=32'h0;
reg	[15:0]	syncEnable_u119_u0=16'h0;
reg	[15:0]	syncEnable_u120_u0=16'h0;
reg		reg_62957a34_u0=1'h0;
wire	[31:0]	mux_u124_u0;
wire		or_u395_u0;
reg		reg_2e3a6914_u0=1'h0;
assign add={31'b0, port_3b9b03c5_}+32'h0;
assign and_u1481_u0=reg_2e3a6914_u0&port_53886836_;
assign subtract={8'b0, port_3b9b03c5_}-9'h1;
assign greaterThanEqualTo_a_signed={subtract[2], subtract[2], subtract[2], subtract[2], subtract[2], subtract[2], subtract[2:0]};
assign greaterThanEqualTo_b_signed=9'h0;
assign greaterThanEqualTo=greaterThanEqualTo_a_signed>=greaterThanEqualTo_b_signed;
assign and_u1482_u0=GO&not_u283_u0;
assign and_u1483_u0=GO&greaterThanEqualTo;
assign not_u283_u0=~greaterThanEqualTo;
assign subtract_u10={8'b0, port_3b9b03c5_}-9'h1;
assign and_u1484_u0=and_u1482_u0&GO;
assign and_u1485_u0=and_u1483_u0&GO;
assign mux_u123=(and_u1484_u0)?9'h2:{subtract_u10[2], subtract_u10[2], subtract_u10[2], subtract_u10[2], subtract_u10[2], subtract_u10[2], subtract_u10[2:0]};
assign add_u47={mux_u123[2], mux_u123[2], mux_u123[2], mux_u123[2], mux_u123[2], mux_u123[2], mux_u123[2], mux_u123[2], mux_u123[2], mux_u123[2], mux_u123[2], mux_u123[2], mux_u123[2], mux_u123[2], mux_u123[2], mux_u123[2], mux_u123[2], mux_u123[2], mux_u123[2], mux_u123[2], mux_u123[2], mux_u123[2], mux_u123[2], mux_u123[2], mux_u123[2], mux_u123[2], mux_u123[2], mux_u123[2], mux_u123[2], mux_u123[2:0]}+32'h0;
assign and_u1486_u0=reg_2e3a6914_u0&port_2d39d825_;
assign and_u1488_u0=reg_62957a34_u0&port_53886836_;
assign add_u48={syncEnable_u119_u0[15], syncEnable_u119_u0}+{port_63c1f3c3_[15], port_63c1f3c3_};
assign subtract_u11=syncEnable_u120_u0-add_u48[16:1];
assign simplePinWrite=16'h1&{16{1'h1}};
assign simplePinWrite_u253=reg_62957a34_u0&{1{reg_62957a34_u0}};
assign simplePinWrite_u254=subtract_u11&{16{reg_62957a34_u0}};
assign simplePinWrite_u255=subtract_u11&{16{reg_62957a34_u0}};
assign simplePinWrite_u256=reg_62957a34_u0&{1{reg_62957a34_u0}};
assign simplePinWrite_u257=16'h1&{16{1'h1}};
always @(posedge CLK)
begin
if (GO)
syncEnable_u117<={add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2:0]};
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u118_u0<=add_u47;
end
always @(posedge CLK)
begin
if (reg_2e3a6914_u0)
syncEnable_u119_u0<=port_768c8415_;
end
always @(posedge CLK)
begin
if (reg_2e3a6914_u0)
syncEnable_u120_u0<=port_63c1f3c3_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_62957a34_u0<=1'h0;
else reg_62957a34_u0<=reg_2e3a6914_u0;
end
assign mux_u124_u0=(reg_2e3a6914_u0)?syncEnable_u117:32'h0;
assign or_u395_u0=reg_2e3a6914_u0|reg_62957a34_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2e3a6914_u0<=1'h0;
else reg_2e3a6914_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u903=1'h0;
assign RESULT_u904=or_u395_u0;
assign RESULT_u905=mux_u124_u0;
assign RESULT_u906=3'h1;
assign RESULT_u907=reg_2e3a6914_u0;
assign RESULT_u908=syncEnable_u118_u0;
assign RESULT_u909=3'h1;
assign RESULT_u910=simplePinWrite_u255;
assign RESULT_u911=simplePinWrite_u253;
assign RESULT_u912=simplePinWrite_u254;
assign RESULT_u913=simplePinWrite;
assign RESULT_u914=simplePinWrite_u257;
assign RESULT_u915=simplePinWrite_u256;
assign DONE=reg_62957a34_u0;
endmodule



module LL1_iunzip_simplememoryreferee_1c6f7bbb_(bus_46f786f5_, bus_3dd26b70_, bus_31d8e4db_, bus_7604351c_, bus_4e6481ad_, bus_6be83458_, bus_2164d186_, bus_51c5d9cf_, bus_010f6c42_, bus_675cdef9_, bus_6f27dbf2_, bus_7943488e_, bus_5c945c19_, bus_5ef9551e_, bus_358645e2_, bus_361af4ce_, bus_1264fa5e_, bus_009a4c19_, bus_6262936b_, bus_35744436_, bus_1dea0faa_, bus_03be4094_, bus_7d72a327_, bus_3946234b_, bus_47c83720_, bus_69d09001_, bus_23f0e20f_, bus_7abd2454_, bus_0ace3741_);
input		bus_46f786f5_;
input		bus_3dd26b70_;
input		bus_31d8e4db_;
input	[15:0]	bus_7604351c_;
input		bus_4e6481ad_;
input	[31:0]	bus_6be83458_;
input	[2:0]	bus_2164d186_;
input		bus_51c5d9cf_;
input	[31:0]	bus_010f6c42_;
input	[2:0]	bus_675cdef9_;
input		bus_6f27dbf2_;
input	[31:0]	bus_7943488e_;
input	[2:0]	bus_5c945c19_;
input		bus_5ef9551e_;
input	[31:0]	bus_358645e2_;
input	[2:0]	bus_361af4ce_;
output	[15:0]	bus_1264fa5e_;
output	[31:0]	bus_009a4c19_;
output		bus_6262936b_;
output		bus_35744436_;
output	[2:0]	bus_1dea0faa_;
output	[15:0]	bus_03be4094_;
output		bus_7d72a327_;
output	[15:0]	bus_3946234b_;
output		bus_47c83720_;
output	[15:0]	bus_69d09001_;
output		bus_23f0e20f_;
output	[15:0]	bus_7abd2454_;
output		bus_0ace3741_;
reg		done_qual_u60_u0=1'h0;
reg		done_qual_u61_u0=1'h0;
reg		done_qual_u62_u0=1'h0;
wire		not_73cf4848_u0;
wire		or_0df849f2_u0;
wire		and_11d4ec5e_u0;
wire		or_620cdf5c_u0;
wire		not_17d4ccc6_u0;
wire		or_20439691_u0;
wire		or_0fa8b73b_u0;
wire		and_11b8746b_u0;
reg		done_qual_u63_u0=1'h0;
wire	[31:0]	mux_2c4fbaa2_u0;
wire		and_73dfd171_u0;
wire		and_44610812_u0;
wire		not_29c81830_u0;
wire		not_006e2a14_u0;
wire		or_5a63991e_u0;
always @(posedge bus_46f786f5_)
begin
if (bus_3dd26b70_)
done_qual_u60_u0<=1'h0;
else done_qual_u60_u0<=bus_5ef9551e_;
end
always @(posedge bus_46f786f5_)
begin
if (bus_3dd26b70_)
done_qual_u61_u0<=1'h0;
else done_qual_u61_u0<=bus_51c5d9cf_;
end
always @(posedge bus_46f786f5_)
begin
if (bus_3dd26b70_)
done_qual_u62_u0<=1'h0;
else done_qual_u62_u0<=bus_4e6481ad_;
end
assign not_73cf4848_u0=~bus_31d8e4db_;
assign or_0df849f2_u0=bus_4e6481ad_|done_qual_u62_u0;
assign and_11d4ec5e_u0=or_0df849f2_u0&bus_31d8e4db_;
assign or_620cdf5c_u0=bus_5ef9551e_|done_qual_u60_u0;
assign not_17d4ccc6_u0=~bus_31d8e4db_;
assign or_20439691_u0=bus_6f27dbf2_|done_qual_u63_u0;
assign or_0fa8b73b_u0=bus_51c5d9cf_|done_qual_u61_u0;
assign and_11b8746b_u0=or_620cdf5c_u0&bus_31d8e4db_;
always @(posedge bus_46f786f5_)
begin
if (bus_3dd26b70_)
done_qual_u63_u0<=1'h0;
else done_qual_u63_u0<=bus_6f27dbf2_;
end
assign mux_2c4fbaa2_u0=({32{bus_4e6481ad_}}&bus_6be83458_)|({32{bus_51c5d9cf_}}&bus_010f6c42_)|({32{bus_6f27dbf2_}}&bus_7943488e_)|({32{bus_5ef9551e_}}&bus_358645e2_);
assign and_73dfd171_u0=or_0fa8b73b_u0&bus_31d8e4db_;
assign and_44610812_u0=or_20439691_u0&bus_31d8e4db_;
assign bus_1264fa5e_=16'h0;
assign bus_009a4c19_=mux_2c4fbaa2_u0;
assign bus_6262936b_=1'h0;
assign bus_35744436_=or_5a63991e_u0;
assign bus_1dea0faa_=3'h1;
assign bus_03be4094_=bus_7604351c_;
assign bus_7d72a327_=and_11d4ec5e_u0;
assign bus_3946234b_=bus_7604351c_;
assign bus_47c83720_=and_73dfd171_u0;
assign bus_69d09001_=bus_7604351c_;
assign bus_23f0e20f_=and_44610812_u0;
assign bus_7abd2454_=bus_7604351c_;
assign bus_0ace3741_=and_11b8746b_u0;
assign not_29c81830_u0=~bus_31d8e4db_;
assign not_006e2a14_u0=~bus_31d8e4db_;
assign or_5a63991e_u0=bus_4e6481ad_|bus_51c5d9cf_|bus_6f27dbf2_|bus_5ef9551e_;
endmodule



module LL1_iunzip_scheduler(CLK, RESET, GO, port_42a101cc_, port_711c21e7_, port_305d8ba1_, port_71394b75_, port_764c2d23_, port_1d25b47a_, port_21a66f1f_, port_7fc5701f_, port_22a38371_, port_31572f8d_, port_411771b7_, port_1b55da6d_, port_10bcdaa8_, port_0379561c_, port_7b10a081_, RESULT, RESULT_u916, RESULT_u917, RESULT_u918, RESULT_u919, RESULT_u920, RESULT_u921, RESULT_u922, RESULT_u923, RESULT_u924, RESULT_u925, RESULT_u926, RESULT_u927, RESULT_u928, RESULT_u929, RESULT_u930, RESULT_u931, RESULT_u932, RESULT_u933, RESULT_u934, DONE);
input		CLK;
input		RESET;
input		GO;
input	[1:0]	port_42a101cc_;
input	[1:0]	port_711c21e7_;
input	[31:0]	port_305d8ba1_;
input	[31:0]	port_71394b75_;
input	[31:0]	port_764c2d23_;
input		port_1d25b47a_;
input		port_21a66f1f_;
input		port_7fc5701f_;
input		port_22a38371_;
input		port_31572f8d_;
input		port_411771b7_;
input		port_1b55da6d_;
input		port_10bcdaa8_;
input		port_0379561c_;
input	[15:0]	port_7b10a081_;
output		RESULT;
output	[1:0]	RESULT_u916;
output		RESULT_u917;
output	[1:0]	RESULT_u918;
output		RESULT_u919;
output	[31:0]	RESULT_u920;
output		RESULT_u921;
output	[31:0]	RESULT_u922;
output		RESULT_u923;
output		RESULT_u924;
output		RESULT_u925;
output	[31:0]	RESULT_u926;
output	[15:0]	RESULT_u927;
output	[2:0]	RESULT_u928;
output		RESULT_u929;
output		RESULT_u930;
output		RESULT_u931;
output		RESULT_u932;
output		RESULT_u933;
output		RESULT_u934;
output		DONE;
wire signed	[31:0]	equals_a_signed;
wire signed	[31:0]	equals_b_signed;
wire		equals;
wire signed	[31:0]	equals_u80_b_signed;
wire		equals_u80;
wire signed	[31:0]	equals_u80_a_signed;
wire signed	[31:0]	equals_u81_b_signed;
wire		equals_u81;
wire signed	[31:0]	equals_u81_a_signed;
wire		equals_u82;
wire signed	[31:0]	equals_u82_b_signed;
wire signed	[31:0]	equals_u82_a_signed;
wire		and_u1490_u0;
wire		and_u1491_u0;
wire		not_u284_u0;
wire		not_u285_u0;
wire		and_u1492_u0;
wire		and_u1493_u0;
wire		simplePinWrite;
reg		reg_09383b58_u0=1'h0;
wire		and_u1494_u0;
reg		reg_09383b58_result_delayed_u0=1'h0;
wire		or_u396_u0;
wire		and_u1495_u0;
reg		and_delayed_u88=1'h0;
wire		or_u397_u0;
wire	[1:0]	mux_u125;
reg		reg_09383b58_result_delayed_result_delayed_u0=1'h0;
wire		and_u1496_u0;
reg		reg_44a467a1_u0=1'h0;
wire		and_u1497_u0;
wire		or_u398_u0;
wire signed	[31:0]	equals_u83_b_signed;
wire signed	[31:0]	equals_u83_a_signed;
wire		equals_u83;
wire		and_u1498_u0;
wire		and_u1499_u0;
wire		not_u286_u0;
wire		not_u287_u0;
wire		and_u1500_u0;
wire		and_u1501_u0;
wire		andOp;
wire		and_u1502_u0;
wire		not_u288_u0;
wire		and_u1503_u0;
wire		simplePinWrite_u258;
wire		and_u1504_u0;
wire		and_u1505_u0;
reg		and_delayed_u89_u0=1'h0;
wire		or_u399_u0;
reg		reg_24bf76a9_u0=1'h0;
reg		and_delayed_u90_u0=1'h0;
wire		not_u289_u0;
wire		and_u1506_u0;
wire		and_u1507_u0;
wire		and_u1508_u0;
wire		and_u1509_u0;
wire		not_u290_u0;
wire		simplePinWrite_u259;
wire		and_u1510_u0;
wire		and_u1511_u0;
wire		or_u400_u0;
reg		reg_20ea2643_u0=1'h0;
reg		and_delayed_u91_u0=1'h0;
reg		reg_20ea2643_result_delayed_u0=1'h0;
reg		and_delayed_u92_u0=1'h0;
wire		and_u1512_u0;
wire		or_u401_u0;
wire		or_u402_u0;
wire	[1:0]	mux_u126_u0;
wire		and_u1513_u0;
reg		and_delayed_u93_u0=1'h0;
wire		or_u403_u0;
wire		and_u1514_u0;
wire		or_u404_u0;
wire	[1:0]	mux_u127_u0;
wire		and_u1515_u0;
wire		and_u1516_u0;
reg		and_delayed_u94_u0=1'h0;
wire		and_u1517_u0;
wire		or_u405_u0;
wire		equals_u84;
wire signed	[31:0]	equals_u84_b_signed;
wire signed	[31:0]	equals_u84_a_signed;
wire		not_u291_u0;
wire		and_u1518_u0;
wire		and_u1519_u0;
wire		and_u1520_u0;
wire		not_u292_u0;
wire		and_u1521_u0;
wire		andOp_u109;
wire		not_u293_u0;
wire		and_u1522_u0;
wire		and_u1523_u0;
wire		simplePinWrite_u260;
reg		reg_1a6d7b26_u0=1'h0;
wire		and_u1524_u0;
wire		or_u406_u0;
wire		and_u1525_u0;
reg		and_delayed_u95_u0=1'h0;
reg		and_delayed_u96_u0=1'h0;
wire		and_u1526_u0;
wire		not_u294_u0;
wire		and_u1527_u0;
wire		and_u1528_u0;
wire		and_u1529_u0;
wire		not_u295_u0;
wire		simplePinWrite_u261;
reg		reg_0807f14a_u0=1'h0;
reg		reg_2d0da07d_u0=1'h0;
wire		or_u407_u0;
wire		and_u1530_u0;
reg		reg_001e3e69_u0=1'h0;
reg		reg_2806cf1c_u0=1'h0;
wire		and_u1531_u0;
wire		and_u1532_u0;
wire		or_u408_u0;
wire	[1:0]	mux_u128_u0;
wire		and_u1533_u0;
reg		and_delayed_u97_u0=1'h0;
wire		or_u409_u0;
wire		and_u1534_u0;
wire	[1:0]	mux_u129_u0;
wire		or_u410_u0;
wire		or_u411_u0;
wire		and_u1535_u0;
wire		or_u412_u0;
reg		reg_41371304_u0=1'h0;
wire		and_u1536_u0;
wire		and_u1537_u0;
wire		equals_u85;
wire signed	[31:0]	equals_u85_a_signed;
wire signed	[31:0]	equals_u85_b_signed;
wire		and_u1538_u0;
wire		and_u1539_u0;
wire		not_u296_u0;
wire signed	[31:0]	lessThan_b_signed;
wire signed	[31:0]	lessThan_a_signed;
wire		lessThan;
wire		and_u1540_u0;
wire		and_u1541_u0;
wire		not_u297_u0;
wire		not_u298_u0;
wire		and_u1542_u0;
wire		and_u1543_u0;
wire		simplePinWrite_u262;
wire	[31:0]	add;
wire		and_u1544_u0;
reg		reg_2d9d5e6b_u0=1'h0;
wire		or_u413_u0;
wire	[31:0]	add_u49;
reg	[15:0]	syncEnable_u121=16'h0;
wire		and_u1545_u0;
reg	[15:0]	syncEnable_u122_u0=16'h0;
reg		and_delayed_u98_u0=1'h0;
wire	[15:0]	mux_u130_u0;
wire		and_u1546_u0;
reg		and_delayed_u99_u0=1'h0;
reg	[2:0]	syncEnable_u123_u0=3'h0;
wire		and_u1547_u0;
wire		and_u1548_u0;
reg	[15:0]	syncEnable_u124_u0=16'h0;
wire	[31:0]	mux_u131_u0;
reg		and_delayed_u100_u0=1'h0;
wire	[15:0]	mux_u132_u0;
reg		and_delayed_u101_u0=1'h0;
reg	[31:0]	syncEnable_u125_u0=32'h0;
wire	[31:0]	mux_u133_u0;
reg		reg_0735f0d2_u0=1'h0;
reg	[15:0]	syncEnable_u126_u0=16'h0;
reg	[31:0]	syncEnable_u127_u0=32'h0;
wire		and_u1549_u0;
wire	[15:0]	mux_u134_u0;
wire		and_u1550_u0;
reg		and_delayed_u102_u0=1'h0;
wire	[1:0]	mux_u135_u0;
wire		or_u414_u0;
wire	[31:0]	mux_u136_u0;
wire		or_u415_u0;
wire		or_u416_u0;
wire	[31:0]	mux_u137_u0;
reg		block_GO_delayed_u2=1'h0;
wire	[1:0]	mux_u138_u0;
wire		or_u417_u0;
reg		scoreboard_7219cf80_reg2=1'h0;
wire		scoreboard_7219cf80_resOr0;
wire		scoreboard_7219cf80_resOr1;
reg		scoreboard_7219cf80_reg0=1'h0;
wire		scoreboard_7219cf80_resOr2;
wire		bus_5d28061f_;
reg		scoreboard_7219cf80_reg1=1'h0;
wire		scoreboard_7219cf80_and;
reg	[31:0]	latch_40712a28_reg=32'h0;
wire	[31:0]	latch_40712a28_out;
reg	[15:0]	latch_62fca6a1_reg=16'h0;
wire	[15:0]	latch_62fca6a1_out;
reg	[2:0]	syncEnable_u128_u0=3'h0;
reg		syncEnable_u129_u0=1'h0;
reg		block_GO_delayed_u3_u0=1'h0;
reg		syncEnable_u130_u0=1'h0;
reg	[31:0]	syncEnable_u131_u0=32'h0;
reg	[15:0]	syncEnable_u132_u0=16'h0;
reg		syncEnable_u133_u0=1'h0;
reg		syncEnable_u134_u0=1'h0;
reg		syncEnable_u135_u0=1'h0;
reg	[31:0]	syncEnable_u136_u0=32'h0;
reg		syncEnable_u137_u0=1'h0;
reg	[31:0]	syncEnable_u138_u0=32'h0;
wire		and_u1551_u0;
reg	[31:0]	fbReg_temp_fsmOldState_LL1_iunzip_1_u0=32'h0;
wire	[31:0]	mux_u139_u0;
wire		or_u418_u0;
reg		loopControl_u1=1'h0;
wire	[15:0]	mux_u140_u0;
reg	[15:0]	fbReg_In1Portvalue_u1=16'h0;
reg		syncEnable_u139_u0=1'h0;
wire		or_u419_u0;
wire		mux_u141_u0;
wire	[1:0]	mux_u142_u0;
wire		or_u420_u0;
reg		reg_7ae9f44d_u0=1'h0;
wire		or_u421_u0;
wire	[31:0]	mux_u143_u0;
reg		reg_7ae9f44d_result_delayed_u0=1'h0;
wire	[31:0]	mux_u144_u0;
wire		or_u422_u0;
wire		or_u423_u0;
wire	[1:0]	mux_u145_u0;
assign equals_a_signed=port_764c2d23_;
assign equals_b_signed=32'h10000;
assign equals=equals_a_signed==equals_b_signed;
assign equals_u80_a_signed=port_764c2d23_;
assign equals_u80_b_signed=32'h10000;
assign equals_u80=equals_u80_a_signed==equals_u80_b_signed;
assign equals_u81_a_signed=port_305d8ba1_;
assign equals_u81_b_signed=32'h2;
assign equals_u81=equals_u81_a_signed==equals_u81_b_signed;
assign equals_u82_a_signed={30'b0, syncEnable_u128_u0[1:0]};
assign equals_u82_b_signed=32'h0;
assign equals_u82=equals_u82_a_signed==equals_u82_b_signed;
assign and_u1490_u0=block_GO_delayed_u3_u0&equals_u82;
assign and_u1491_u0=block_GO_delayed_u3_u0&not_u284_u0;
assign not_u284_u0=~equals_u82;
assign not_u285_u0=~syncEnable_u129_u0;
assign and_u1492_u0=and_u1496_u0&not_u285_u0;
assign and_u1493_u0=and_u1496_u0&syncEnable_u129_u0;
assign simplePinWrite=and_u1494_u0&{1{and_u1494_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_09383b58_u0<=1'h0;
else reg_09383b58_u0<=and_u1494_u0;
end
assign and_u1494_u0=and_u1493_u0&and_u1496_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_09383b58_result_delayed_u0<=1'h0;
else reg_09383b58_result_delayed_u0<=reg_09383b58_u0;
end
assign or_u396_u0=reg_09383b58_result_delayed_result_delayed_u0|and_delayed_u88;
assign and_u1495_u0=and_u1492_u0&and_u1496_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u88<=1'h0;
else and_delayed_u88<=and_u1495_u0;
end
assign or_u397_u0=and_u1494_u0|and_u1495_u0;
assign mux_u125=(and_u1494_u0)?2'h1:2'h3;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_09383b58_result_delayed_result_delayed_u0<=1'h0;
else reg_09383b58_result_delayed_result_delayed_u0<=reg_09383b58_result_delayed_u0;
end
assign and_u1496_u0=and_u1490_u0&block_GO_delayed_u3_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_44a467a1_u0<=1'h0;
else reg_44a467a1_u0<=and_u1497_u0;
end
assign and_u1497_u0=and_u1491_u0&block_GO_delayed_u3_u0;
assign or_u398_u0=or_u396_u0|reg_44a467a1_u0;
assign equals_u83_a_signed={30'b0, syncEnable_u128_u0[1:0]};
assign equals_u83_b_signed=32'h1;
assign equals_u83=equals_u83_a_signed==equals_u83_b_signed;
assign and_u1498_u0=block_GO_delayed_u3_u0&equals_u83;
assign and_u1499_u0=block_GO_delayed_u3_u0&not_u286_u0;
assign not_u286_u0=~equals_u83;
assign not_u287_u0=~syncEnable_u133_u0;
assign and_u1500_u0=and_u1517_u0&syncEnable_u133_u0;
assign and_u1501_u0=and_u1517_u0&not_u287_u0;
assign andOp=port_22a38371_&port_31572f8d_;
assign and_u1502_u0=and_u1514_u0&not_u288_u0;
assign not_u288_u0=~andOp;
assign and_u1503_u0=and_u1514_u0&andOp;
assign simplePinWrite_u258=and_u1505_u0&{1{and_u1505_u0}};
assign and_u1504_u0=and_u1502_u0&and_u1514_u0;
assign and_u1505_u0=and_u1503_u0&and_u1514_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u89_u0<=1'h0;
else and_delayed_u89_u0<=and_u1504_u0;
end
assign or_u399_u0=and_delayed_u89_u0|reg_24bf76a9_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_24bf76a9_u0<=1'h0;
else reg_24bf76a9_u0<=and_delayed_u90_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u90_u0<=1'h0;
else and_delayed_u90_u0<=and_u1505_u0;
end
assign not_u289_u0=~syncEnable_u130_u0;
assign and_u1506_u0=and_u1515_u0&not_u289_u0;
assign and_u1507_u0=and_u1515_u0&syncEnable_u130_u0;
assign and_u1508_u0=and_u1513_u0&port_22a38371_;
assign and_u1509_u0=and_u1513_u0&not_u290_u0;
assign not_u290_u0=~port_22a38371_;
assign simplePinWrite_u259=and_u1511_u0&{1{and_u1511_u0}};
assign and_u1510_u0=and_u1509_u0&and_u1513_u0;
assign and_u1511_u0=and_u1508_u0&and_u1513_u0;
assign or_u400_u0=and_delayed_u92_u0|reg_20ea2643_result_delayed_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_20ea2643_u0<=1'h0;
else reg_20ea2643_u0<=and_delayed_u91_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u91_u0<=1'h0;
else and_delayed_u91_u0<=and_u1511_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_20ea2643_result_delayed_u0<=1'h0;
else reg_20ea2643_result_delayed_u0<=reg_20ea2643_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u92_u0<=1'h0;
else and_delayed_u92_u0<=and_u1510_u0;
end
assign and_u1512_u0=and_u1506_u0&and_u1515_u0;
assign or_u401_u0=or_u400_u0|and_delayed_u93_u0;
assign or_u402_u0=and_u1511_u0|and_u1512_u0;
assign mux_u126_u0=(and_u1511_u0)?2'h2:2'h3;
assign and_u1513_u0=and_u1507_u0&and_u1515_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u93_u0<=1'h0;
else and_delayed_u93_u0<=and_u1512_u0;
end
assign or_u403_u0=or_u399_u0|or_u401_u0;
assign and_u1514_u0=and_u1500_u0&and_u1517_u0;
assign or_u404_u0=and_u1505_u0|or_u402_u0;
assign mux_u127_u0=(and_u1505_u0)?2'h0:{1'b1, mux_u126_u0[0]};
assign and_u1515_u0=and_u1501_u0&and_u1517_u0;
assign and_u1516_u0=and_u1499_u0&block_GO_delayed_u3_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u94_u0<=1'h0;
else and_delayed_u94_u0<=and_u1516_u0;
end
assign and_u1517_u0=and_u1498_u0&block_GO_delayed_u3_u0;
assign or_u405_u0=or_u403_u0|and_delayed_u94_u0;
assign equals_u84_a_signed={30'b0, syncEnable_u128_u0[1:0]};
assign equals_u84_b_signed=32'h2;
assign equals_u84=equals_u84_a_signed==equals_u84_b_signed;
assign not_u291_u0=~equals_u84;
assign and_u1518_u0=block_GO_delayed_u3_u0&equals_u84;
assign and_u1519_u0=block_GO_delayed_u3_u0&not_u291_u0;
assign and_u1520_u0=and_u1537_u0&not_u292_u0;
assign not_u292_u0=~syncEnable_u135_u0;
assign and_u1521_u0=and_u1537_u0&syncEnable_u135_u0;
assign andOp_u109=port_22a38371_&port_31572f8d_;
assign not_u293_u0=~andOp_u109;
assign and_u1522_u0=and_u1535_u0&not_u293_u0;
assign and_u1523_u0=and_u1535_u0&andOp_u109;
assign simplePinWrite_u260=and_u1525_u0&{1{and_u1525_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1a6d7b26_u0<=1'h0;
else reg_1a6d7b26_u0<=and_delayed_u96_u0;
end
assign and_u1524_u0=and_u1522_u0&and_u1535_u0;
assign or_u406_u0=and_delayed_u95_u0|reg_1a6d7b26_u0;
assign and_u1525_u0=and_u1523_u0&and_u1535_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u95_u0<=1'h0;
else and_delayed_u95_u0<=and_u1524_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u96_u0<=1'h0;
else and_delayed_u96_u0<=and_u1525_u0;
end
assign and_u1526_u0=and_u1534_u0&syncEnable_u134_u0;
assign not_u294_u0=~syncEnable_u134_u0;
assign and_u1527_u0=and_u1534_u0&not_u294_u0;
assign and_u1528_u0=and_u1533_u0&not_u295_u0;
assign and_u1529_u0=and_u1533_u0&port_31572f8d_;
assign not_u295_u0=~port_31572f8d_;
assign simplePinWrite_u261=and_u1531_u0&{1{and_u1531_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0807f14a_u0<=1'h0;
else reg_0807f14a_u0<=reg_001e3e69_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2d0da07d_u0<=1'h0;
else reg_2d0da07d_u0<=and_u1530_u0;
end
assign or_u407_u0=reg_0807f14a_u0|reg_2d0da07d_u0;
assign and_u1530_u0=and_u1528_u0&and_u1533_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_001e3e69_u0<=1'h0;
else reg_001e3e69_u0<=reg_2806cf1c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2806cf1c_u0<=1'h0;
else reg_2806cf1c_u0<=and_u1531_u0;
end
assign and_u1531_u0=and_u1529_u0&and_u1533_u0;
assign and_u1532_u0=and_u1527_u0&and_u1534_u0;
assign or_u408_u0=and_u1531_u0|and_u1532_u0;
assign mux_u128_u0=(and_u1531_u0)?2'h1:2'h3;
assign and_u1533_u0=and_u1526_u0&and_u1534_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u97_u0<=1'h0;
else and_delayed_u97_u0<=and_u1532_u0;
end
assign or_u409_u0=or_u407_u0|and_delayed_u97_u0;
assign and_u1534_u0=and_u1520_u0&and_u1537_u0;
assign mux_u129_u0=(and_u1525_u0)?2'h0:{mux_u128_u0[1], 1'b1};
assign or_u410_u0=and_u1525_u0|or_u408_u0;
assign or_u411_u0=or_u406_u0|or_u409_u0;
assign and_u1535_u0=and_u1521_u0&and_u1537_u0;
assign or_u412_u0=reg_41371304_u0|or_u411_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_41371304_u0<=1'h0;
else reg_41371304_u0<=and_u1536_u0;
end
assign and_u1536_u0=and_u1519_u0&block_GO_delayed_u3_u0;
assign and_u1537_u0=and_u1518_u0&block_GO_delayed_u3_u0;
assign equals_u85_a_signed={30'b0, syncEnable_u128_u0[1:0]};
assign equals_u85_b_signed=32'h3;
assign equals_u85=equals_u85_a_signed==equals_u85_b_signed;
assign and_u1538_u0=block_GO_delayed_u3_u0&equals_u85;
assign and_u1539_u0=block_GO_delayed_u3_u0&not_u296_u0;
assign not_u296_u0=~equals_u85;
assign lessThan_a_signed=syncEnable_u138_u0;
assign lessThan_b_signed=syncEnable_u136_u0;
assign lessThan=lessThan_a_signed<lessThan_b_signed;
assign and_u1540_u0=and_u1549_u0&lessThan;
assign and_u1541_u0=and_u1549_u0&not_u297_u0;
assign not_u297_u0=~lessThan;
assign not_u298_u0=~syncEnable_u137_u0;
assign and_u1542_u0=and_u1548_u0&not_u298_u0;
assign and_u1543_u0=and_u1548_u0&syncEnable_u137_u0;
assign simplePinWrite_u262=and_u1545_u0&{1{and_u1545_u0}};
assign add=syncEnable_u138_u0+32'h0;
assign and_u1544_u0=reg_2d9d5e6b_u0&port_1d25b47a_;
always @(posedge CLK or posedge and_u1545_u0 or posedge or_u413_u0)
begin
if (or_u413_u0)
reg_2d9d5e6b_u0<=1'h0;
else if (and_u1545_u0)
reg_2d9d5e6b_u0<=1'h1;
else reg_2d9d5e6b_u0<=reg_2d9d5e6b_u0;
end
assign or_u413_u0=and_u1544_u0|RESET;
assign add_u49=syncEnable_u138_u0+32'h1;
always @(posedge CLK)
begin
if (and_u1545_u0)
syncEnable_u121<=port_7b10a081_;
end
assign and_u1545_u0=and_u1543_u0&and_u1548_u0;
always @(posedge CLK)
begin
if (and_u1548_u0)
syncEnable_u122_u0<=syncEnable_u132_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u98_u0<=1'h0;
else and_delayed_u98_u0<=and_u1545_u0;
end
assign mux_u130_u0=(and_delayed_u98_u0)?syncEnable_u121:syncEnable_u122_u0;
assign and_u1546_u0=and_u1542_u0&and_u1548_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u99_u0<=1'h0;
else and_delayed_u99_u0<=and_u1546_u0;
end
always @(posedge CLK)
begin
if (and_u1547_u0)
syncEnable_u123_u0<={1'b0, port_42a101cc_};
end
assign and_u1547_u0=and_u1541_u0&and_u1549_u0;
assign and_u1548_u0=and_u1540_u0&and_u1549_u0;
always @(posedge CLK)
begin
if (and_u1549_u0)
syncEnable_u124_u0<=syncEnable_u132_u0;
end
assign mux_u131_u0=(and_delayed_u101_u0)?syncEnable_u125_u0:{30'b0, syncEnable_u123_u0[1:0]};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u100_u0<=1'h0;
else and_delayed_u100_u0<=and_u1547_u0;
end
assign mux_u132_u0=(and_delayed_u101_u0)?mux_u130_u0:syncEnable_u124_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u101_u0<=1'h0;
else and_delayed_u101_u0<=and_u1548_u0;
end
always @(posedge CLK)
begin
if (and_u1549_u0)
syncEnable_u125_u0<=syncEnable_u131_u0;
end
assign mux_u133_u0=(reg_0735f0d2_u0)?mux_u131_u0:syncEnable_u127_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0735f0d2_u0<=1'h0;
else reg_0735f0d2_u0<=and_u1549_u0;
end
always @(posedge CLK)
begin
if (block_GO_delayed_u3_u0)
syncEnable_u126_u0<=syncEnable_u132_u0;
end
always @(posedge CLK)
begin
if (block_GO_delayed_u3_u0)
syncEnable_u127_u0<=syncEnable_u131_u0;
end
assign and_u1549_u0=and_u1538_u0&block_GO_delayed_u3_u0;
assign mux_u134_u0=(reg_0735f0d2_u0)?mux_u132_u0:syncEnable_u126_u0;
assign and_u1550_u0=and_u1539_u0&block_GO_delayed_u3_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u102_u0<=1'h0;
else and_delayed_u102_u0<=and_u1550_u0;
end
assign mux_u135_u0=({2{or_u397_u0}}&{mux_u125[1], 1'b1})|({2{or_u404_u0}}&mux_u127_u0)|({2{or_u410_u0}}&mux_u129_u0)|({2{and_u1547_u0}}&port_42a101cc_);
assign or_u414_u0=or_u397_u0|or_u404_u0|or_u410_u0|and_u1547_u0;
assign mux_u136_u0=(and_u1495_u0)?32'h0:32'hfffffffd;
assign or_u415_u0=and_u1495_u0|and_u1547_u0;
assign or_u416_u0=and_u1494_u0|and_u1545_u0;
assign mux_u137_u0=(and_u1494_u0)?32'h0:add_u49;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
block_GO_delayed_u2<=1'h0;
else block_GO_delayed_u2<=block_GO_delayed_u3_u0;
end
assign mux_u138_u0=({2{and_u1495_u0}}&2'h0)|({2{and_u1512_u0}}&2'h1)|({2{and_u1532_u0}}&2'h2);
assign or_u417_u0=and_u1495_u0|and_u1512_u0|and_u1532_u0;
always @(posedge CLK)
begin
if (bus_5d28061f_)
scoreboard_7219cf80_reg2<=1'h0;
else if (or_u405_u0)
scoreboard_7219cf80_reg2<=1'h1;
else scoreboard_7219cf80_reg2<=scoreboard_7219cf80_reg2;
end
assign scoreboard_7219cf80_resOr0=or_u412_u0|scoreboard_7219cf80_reg0;
assign scoreboard_7219cf80_resOr1=or_u398_u0|scoreboard_7219cf80_reg1;
always @(posedge CLK)
begin
if (bus_5d28061f_)
scoreboard_7219cf80_reg0<=1'h0;
else if (or_u412_u0)
scoreboard_7219cf80_reg0<=1'h1;
else scoreboard_7219cf80_reg0<=scoreboard_7219cf80_reg0;
end
assign scoreboard_7219cf80_resOr2=or_u405_u0|scoreboard_7219cf80_reg2;
assign bus_5d28061f_=scoreboard_7219cf80_and|RESET;
always @(posedge CLK)
begin
if (bus_5d28061f_)
scoreboard_7219cf80_reg1<=1'h0;
else if (or_u398_u0)
scoreboard_7219cf80_reg1<=1'h1;
else scoreboard_7219cf80_reg1<=scoreboard_7219cf80_reg1;
end
assign scoreboard_7219cf80_and=scoreboard_7219cf80_resOr0&scoreboard_7219cf80_resOr1&scoreboard_7219cf80_resOr2;
always @(posedge CLK)
begin
if (block_GO_delayed_u2)
latch_40712a28_reg<=mux_u133_u0;
end
assign latch_40712a28_out=(block_GO_delayed_u2)?mux_u133_u0:latch_40712a28_reg;
always @(posedge CLK)
begin
if (block_GO_delayed_u2)
latch_62fca6a1_reg<=mux_u134_u0;
end
assign latch_62fca6a1_out=(block_GO_delayed_u2)?mux_u134_u0:latch_62fca6a1_reg;
always @(posedge CLK)
begin
if (and_u1551_u0)
syncEnable_u128_u0<={1'b0, port_711c21e7_};
end
always @(posedge CLK)
begin
if (and_u1551_u0)
syncEnable_u129_u0<=equals_u81;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
block_GO_delayed_u3_u0<=1'h0;
else block_GO_delayed_u3_u0<=and_u1551_u0;
end
always @(posedge CLK)
begin
if (and_u1551_u0)
syncEnable_u130_u0<=port_21a66f1f_;
end
always @(posedge CLK)
begin
if (and_u1551_u0)
syncEnable_u131_u0<=mux_u139_u0;
end
always @(posedge CLK)
begin
if (and_u1551_u0)
syncEnable_u132_u0<=mux_u140_u0;
end
always @(posedge CLK)
begin
if (and_u1551_u0)
syncEnable_u133_u0<=equals;
end
always @(posedge CLK)
begin
if (and_u1551_u0)
syncEnable_u134_u0<=port_21a66f1f_;
end
always @(posedge CLK)
begin
if (and_u1551_u0)
syncEnable_u135_u0<=equals_u80;
end
always @(posedge CLK)
begin
if (and_u1551_u0)
syncEnable_u136_u0<=port_71394b75_;
end
always @(posedge CLK)
begin
if (and_u1551_u0)
syncEnable_u137_u0<=port_21a66f1f_;
end
always @(posedge CLK)
begin
if (and_u1551_u0)
syncEnable_u138_u0<=port_305d8ba1_;
end
assign and_u1551_u0=or_u418_u0&or_u418_u0;
always @(posedge CLK)
begin
if (scoreboard_7219cf80_and)
fbReg_temp_fsmOldState_LL1_iunzip_1_u0<=latch_40712a28_out;
end
assign mux_u139_u0=(reg_7ae9f44d_result_delayed_u0)?32'h0:fbReg_temp_fsmOldState_LL1_iunzip_1_u0;
assign or_u418_u0=reg_7ae9f44d_result_delayed_u0|loopControl_u1;
always @(posedge CLK or posedge syncEnable_u139_u0)
begin
if (syncEnable_u139_u0)
loopControl_u1<=1'h0;
else loopControl_u1<=scoreboard_7219cf80_and;
end
assign mux_u140_u0=(reg_7ae9f44d_result_delayed_u0)?16'h0:fbReg_In1Portvalue_u1;
always @(posedge CLK)
begin
if (scoreboard_7219cf80_and)
fbReg_In1Portvalue_u1<=latch_62fca6a1_out;
end
always @(posedge CLK)
begin
if (reg_7ae9f44d_result_delayed_u0)
syncEnable_u139_u0<=RESET;
end
assign or_u419_u0=GO|and_u1495_u0;
assign mux_u141_u0=(GO)?1'h0:1'h1;
assign mux_u142_u0=(GO)?2'h0:mux_u138_u0;
assign or_u420_u0=GO|or_u417_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7ae9f44d_u0<=1'h0;
else reg_7ae9f44d_u0<=GO;
end
assign or_u421_u0=GO|or_u416_u0;
assign mux_u143_u0=(GO)?32'h0:mux_u137_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7ae9f44d_result_delayed_u0<=1'h0;
else reg_7ae9f44d_result_delayed_u0<=reg_7ae9f44d_u0;
end
assign mux_u144_u0=(GO)?32'hfffffffd:{mux_u136_u0[31:2], 1'b0, mux_u136_u0[0]};
assign or_u422_u0=GO|or_u415_u0;
assign or_u423_u0=GO|or_u414_u0;
assign mux_u145_u0=(GO)?2'h0:mux_u135_u0;
assign RESULT=or_u420_u0;
assign RESULT_u916=mux_u142_u0;
assign RESULT_u917=or_u423_u0;
assign RESULT_u918=mux_u145_u0;
assign RESULT_u919=or_u421_u0;
assign RESULT_u920=mux_u143_u0;
assign RESULT_u921=or_u422_u0;
assign RESULT_u922={mux_u144_u0[31:2], 1'b0, mux_u144_u0[0]};
assign RESULT_u923=or_u419_u0;
assign RESULT_u924=mux_u141_u0;
assign RESULT_u925=and_u1545_u0;
assign RESULT_u926=add;
assign RESULT_u927=port_7b10a081_;
assign RESULT_u928=3'h1;
assign RESULT_u929=simplePinWrite_u262;
assign RESULT_u930=simplePinWrite_u259;
assign RESULT_u931=simplePinWrite_u258;
assign RESULT_u932=simplePinWrite_u260;
assign RESULT_u933=simplePinWrite_u261;
assign RESULT_u934=simplePinWrite;
assign DONE=1'h0;
endmodule



module LL1_iunzip_globalreset_physical_7bb59c58_(bus_0bf03daf_, bus_7876706a_, bus_1a0482e7_);
input		bus_0bf03daf_;
input		bus_7876706a_;
output		bus_1a0482e7_;
reg		sample_u22=1'h0;
wire		not_413c03fc_u0;
wire		or_3dcc81fd_u0;
reg		cross_u22=1'h0;
wire		and_47e34a17_u0;
reg		final_u22=1'h1;
reg		glitch_u22=1'h0;
always @(posedge bus_0bf03daf_)
begin
sample_u22<=1'h1;
end
assign not_413c03fc_u0=~and_47e34a17_u0;
assign or_3dcc81fd_u0=bus_7876706a_|final_u22;
assign bus_1a0482e7_=or_3dcc81fd_u0;
always @(posedge bus_0bf03daf_)
begin
cross_u22<=sample_u22;
end
assign and_47e34a17_u0=cross_u22&glitch_u22;
always @(posedge bus_0bf03daf_)
begin
final_u22<=not_413c03fc_u0;
end
always @(posedge bus_0bf03daf_)
begin
glitch_u22<=cross_u22;
end
endmodule


