// __  ___ __ ___  _ __   ___  ___ 
// \ \/ / '__/ _ \| '_ \ / _ \/ __|
//  >  <| | | (_) | | | | (_) \__ \
// /_/\_\_|  \___/|_| |_|\___/|___/
// 
// Xronos synthesizer version
// Run date: Thu 2 Nov 2017 13:59:19 +0000
// 

module resized_LH1_xy(In1_ACK, Out1_ACK, Out1_DATA, In1_SEND, Out1_RDY, CLK, In1_DATA, In1_COUNT, Out1_COUNT, RESET, Out1_SEND);
wire		consumeRow_go;
output		In1_ACK;
input		Out1_ACK;
wire		consumeRow_done;
output	[15:0]	Out1_DATA;
input		In1_SEND;
input		Out1_RDY;
input		CLK;
input	[15:0]	In1_DATA;
wire		reset_done;
wire		repeatRowExpanded_go;
wire		reset_go;
input	[15:0]	In1_COUNT;
output	[15:0]	Out1_COUNT;
input		RESET;
output		Out1_SEND;
wire		repeatRowExpanded_done;
wire		bus_146eb89f_;
wire		bus_0fe08b68_;
wire	[15:0]	bus_37dd7726_;
wire		bus_2698717b_;
wire	[15:0]	bus_72d7955d_;
wire		bus_67d19bcd_;
wire	[31:0]	bus_3d2b1c2b_;
wire		bus_71c557ad_;
wire		bus_2d657228_;
wire	[15:0]	reset_u9;
wire		reset_u10;
wire		resized_LH1_xy_reset_instance_DONE;
wire		reset;
wire	[15:0]	reset_u11;
wire		bus_1823b71b_;
wire	[31:0]	bus_0dea0337_;
wire		bus_053c348c_;
wire		bus_41a72575_;
wire	[15:0]	bus_043f5796_;
wire		bus_47674f00_;
wire	[2:0]	bus_54d5acc6_;
wire	[15:0]	bus_5d969c8b_;
wire		bus_4a047406_;
wire		bus_382ad4dd_;
wire		repeatRowExpanded_u28;
wire	[2:0]	repeatRowExpanded_u31;
wire		repeatRowExpanded;
wire	[15:0]	repeatRowExpanded_u24;
wire	[15:0]	repeatRowExpanded_u30;
wire		resized_LH1_xy_repeatRowExpanded_instance_DONE;
wire		repeatRowExpanded_u25;
wire	[2:0]	repeatRowExpanded_u27;
wire	[31:0]	repeatRowExpanded_u29;
wire	[31:0]	repeatRowExpanded_u26;
wire	[2:0]	bus_527ad470_;
wire		bus_7cc52ea4_;
wire		bus_6818c058_;
wire	[15:0]	bus_17060ee9_;
wire		bus_7232d2ee_;
wire	[31:0]	bus_1c368516_;
wire		bus_44b70675_;
wire	[15:0]	bus_0af0ab39_;
wire		bus_178082e9_;
wire		scheduler_u267;
wire		scheduler_u281;
wire	[31:0]	scheduler_u272;
wire		resized_LH1_xy_scheduler_instance_DONE;
wire		scheduler_u275;
wire	[31:0]	scheduler_u266;
wire	[2:0]	scheduler_u277;
wire		scheduler;
wire		scheduler_u269;
wire	[31:0]	scheduler_u270;
wire		scheduler_u283;
wire		scheduler_u273;
wire		scheduler_u280;
wire		scheduler_u271;
wire	[15:0]	scheduler_u279;
wire		scheduler_u278;
wire	[15:0]	scheduler_u282;
wire		scheduler_u274;
wire	[31:0]	scheduler_u276;
wire		scheduler_u268;
wire	[31:0]	bus_4a96edb8_;
wire	[31:0]	bus_7668b64d_;
wire	[15:0]	bus_70ada90a_;
wire	[15:0]	bus_2d676b21_;
wire		bus_6bc2d2f4_;
wire	[15:0]	consumeRow_u30;
wire		consumeRow_u31;
wire	[31:0]	consumeRow_u36;
wire		consumeRow;
wire	[15:0]	consumeRow_u33;
wire	[15:0]	consumeRow_u37;
wire		resized_LH1_xy_consumeRow_instance_DONE;
wire	[31:0]	consumeRow_u32;
wire	[2:0]	consumeRow_u34;
wire		consumeRow_u39;
wire	[2:0]	consumeRow_u38;
wire		consumeRow_u35;
assign consumeRow_go=scheduler_u278;
assign In1_ACK=consumeRow_u39;
assign consumeRow_done=bus_4a047406_;
assign Out1_DATA=scheduler_u282;
assign reset_done=bus_2d657228_;
assign repeatRowExpanded_go=scheduler_u280;
assign reset_go=scheduler_u281;
assign Out1_COUNT=scheduler_u279;
assign Out1_SEND=scheduler_u283;
assign repeatRowExpanded_done=bus_71c557ad_;
resized_LH1_xy_Kicker_43 resized_LH1_xy_Kicker_43_1(.CLK(CLK), .RESET(bus_67d19bcd_), 
  .bus_146eb89f_(bus_146eb89f_));
resized_LH1_xy_structuralmemory_2108298e_ resized_LH1_xy_structuralmemory_2108298e__1(.CLK_u17(CLK), 
  .bus_3a8ce0e8_(bus_67d19bcd_), .bus_32b68420_(bus_0dea0337_), .bus_4efd6486_(3'h1), 
  .bus_677fabb8_(bus_41a72575_), .bus_1c42c4da_(bus_47674f00_), .bus_5d26b9a7_(bus_043f5796_), 
  .bus_37dd7726_(bus_37dd7726_), .bus_0fe08b68_(bus_0fe08b68_));
resized_LH1_xy_stateVar_Out1PortEnable resized_LH1_xy_stateVar_Out1PortEnable_1(.bus_7dadb443_(CLK), 
  .bus_2cfd1fd9_(bus_67d19bcd_), .bus_105e9f86_(scheduler_u273), .bus_4406fa74_(scheduler_u274), 
  .bus_2698717b_(bus_2698717b_));
resized_LH1_xy_stateVar_x resized_LH1_xy_stateVar_x_1(.bus_78bae313_(CLK), .bus_6b0a580d_(bus_67d19bcd_), 
  .bus_4a98ed23_(consumeRow), .bus_5ce6cb87_(consumeRow_u30), .bus_3e718195_(reset_u10), 
  .bus_18105192_(16'h0), .bus_72d7955d_(bus_72d7955d_));
resized_LH1_xy_globalreset_physical_790ef242_ resized_LH1_xy_globalreset_physical_790ef242__1(.bus_664d27ed_(CLK), 
  .bus_42d18000_(RESET), .bus_67d19bcd_(bus_67d19bcd_));
resized_LH1_xy_stateVar_fsmOldState_resized_LH1_xy resized_LH1_xy_stateVar_fsmOldState_resized_LH1_xy_1(.bus_201216da_(CLK), 
  .bus_66f3f92d_(bus_67d19bcd_), .bus_7673123e_(scheduler), .bus_3fa4cd9c_(32'h0), 
  .bus_3d2b1c2b_(bus_3d2b1c2b_));
assign bus_71c557ad_=resized_LH1_xy_repeatRowExpanded_instance_DONE&{1{resized_LH1_xy_repeatRowExpanded_instance_DONE}};
assign bus_2d657228_=resized_LH1_xy_reset_instance_DONE&{1{resized_LH1_xy_reset_instance_DONE}};
resized_LH1_xy_reset resized_LH1_xy_reset_instance(.CLK(CLK), .RESET(bus_67d19bcd_), 
  .GO(reset_go), .DONE(resized_LH1_xy_reset_instance_DONE), .RESULT(reset), .RESULT_u1852(reset_u9), 
  .RESULT_u1853(reset_u10), .RESULT_u1854(reset_u11));
resized_LH1_xy_simplememoryreferee_07b85719_ resized_LH1_xy_simplememoryreferee_07b85719__1(.bus_0b291028_(CLK), 
  .bus_154448d0_(bus_67d19bcd_), .bus_2afbec8d_(bus_0fe08b68_), .bus_1f157a32_(bus_37dd7726_), 
  .bus_6d609752_(consumeRow_u35), .bus_5486e989_(consumeRow_u37), .bus_25b9b8db_(consumeRow_u36), 
  .bus_0756d9ea_(3'h1), .bus_588863ee_(repeatRowExpanded_u25), .bus_79191f33_(repeatRowExpanded_u26), 
  .bus_4bdb631c_(3'h1), .bus_043f5796_(bus_043f5796_), .bus_0dea0337_(bus_0dea0337_), 
  .bus_47674f00_(bus_47674f00_), .bus_41a72575_(bus_41a72575_), .bus_54d5acc6_(bus_54d5acc6_), 
  .bus_1823b71b_(bus_1823b71b_), .bus_5d969c8b_(bus_5d969c8b_), .bus_053c348c_(bus_053c348c_));
assign bus_4a047406_=resized_LH1_xy_consumeRow_instance_DONE&{1{resized_LH1_xy_consumeRow_instance_DONE}};
resized_LH1_xy_stateVar_fsmState_resized_LH1_xy resized_LH1_xy_stateVar_fsmState_resized_LH1_xy_1(.bus_3631bc0b_(CLK), 
  .bus_0708d8fb_(bus_67d19bcd_), .bus_4602c2a7_(scheduler_u267), .bus_3c662fde_(scheduler_u268), 
  .bus_382ad4dd_(bus_382ad4dd_));
resized_LH1_xy_repeatRowExpanded resized_LH1_xy_repeatRowExpanded_instance(.CLK(CLK), 
  .RESET(bus_67d19bcd_), .GO(repeatRowExpanded_go), .port_1819de90_(bus_70ada90a_), 
  .port_5d43c181_(bus_053c348c_), .port_00ba0d3b_(bus_5d969c8b_), .port_6635e8af_(bus_6818c058_), 
  .DONE(resized_LH1_xy_repeatRowExpanded_instance_DONE), .RESULT(repeatRowExpanded), 
  .RESULT_u1855(repeatRowExpanded_u24), .RESULT_u1856(repeatRowExpanded_u25), 
  .RESULT_u1857(repeatRowExpanded_u26), .RESULT_u1858(repeatRowExpanded_u27), 
  .RESULT_u1859(repeatRowExpanded_u28), .RESULT_u1860(repeatRowExpanded_u29), 
  .RESULT_u1861(repeatRowExpanded_u30), .RESULT_u1862(repeatRowExpanded_u31));
resized_LH1_xy_simplememoryreferee_4f8eca27_ resized_LH1_xy_simplememoryreferee_4f8eca27__1(.bus_13a35abe_(CLK), 
  .bus_537d7f21_(bus_67d19bcd_), .bus_67df8591_(bus_6bc2d2f4_), .bus_26c151a5_(bus_2d676b21_), 
  .bus_7e206820_(consumeRow_u31), .bus_0bdb3367_(consumeRow_u33), .bus_3ac51013_(consumeRow_u32), 
  .bus_7de908f2_(3'h1), .bus_2043bfd1_(repeatRowExpanded_u28), .bus_0ca641af_(repeatRowExpanded_u30), 
  .bus_6077dae8_(repeatRowExpanded_u29), .bus_0fd5a0d9_(3'h1), .bus_2444a5e9_(scheduler_u275), 
  .bus_242bf648_(scheduler_u276), .bus_528d16c5_(3'h1), .bus_17060ee9_(bus_17060ee9_), 
  .bus_1c368516_(bus_1c368516_), .bus_178082e9_(bus_178082e9_), .bus_44b70675_(bus_44b70675_), 
  .bus_527ad470_(bus_527ad470_), .bus_7232d2ee_(bus_7232d2ee_), .bus_6818c058_(bus_6818c058_), 
  .bus_0af0ab39_(bus_0af0ab39_), .bus_7cc52ea4_(bus_7cc52ea4_));
resized_LH1_xy_scheduler resized_LH1_xy_scheduler_instance(.CLK(CLK), .RESET(bus_67d19bcd_), 
  .GO(bus_146eb89f_), .port_6105e58c_(32'h0), .port_0a81f2c6_(bus_382ad4dd_), .port_3bb784d0_(bus_4a96edb8_), 
  .port_1ca215c6_(bus_7668b64d_), .port_5071c1a7_(bus_2698717b_), .port_008a440f_(bus_72d7955d_), 
  .port_1ba874b3_(bus_70ada90a_), .port_63d562ec_(bus_7cc52ea4_), .port_2ccab656_(bus_0af0ab39_), 
  .port_2adbeb14_(Out1_RDY), .port_218764d5_(reset_done), .port_51b44ade_(consumeRow_done), 
  .port_58303e5a_(In1_SEND), .port_1be35c61_(repeatRowExpanded_done), .DONE(resized_LH1_xy_scheduler_instance_DONE), 
  .RESULT(scheduler), .RESULT_u1863(scheduler_u266), .RESULT_u1864(scheduler_u267), 
  .RESULT_u1865(scheduler_u268), .RESULT_u1866(scheduler_u269), .RESULT_u1867(scheduler_u270), 
  .RESULT_u1868(scheduler_u271), .RESULT_u1869(scheduler_u272), .RESULT_u1870(scheduler_u273), 
  .RESULT_u1871(scheduler_u274), .RESULT_u1872(scheduler_u275), .RESULT_u1873(scheduler_u276), 
  .RESULT_u1874(scheduler_u277), .RESULT_u1875(scheduler_u278), .RESULT_u1876(scheduler_u279), 
  .RESULT_u1877(scheduler_u280), .RESULT_u1878(scheduler_u281), .RESULT_u1879(scheduler_u282), 
  .RESULT_u1880(scheduler_u283));
resized_LH1_xy_stateVar_Out1TokenIndex resized_LH1_xy_stateVar_Out1TokenIndex_1(.bus_44763466_(CLK), 
  .bus_08eb61b0_(bus_67d19bcd_), .bus_3d7dc20a_(scheduler_u269), .bus_1be81a8d_(scheduler_u270), 
  .bus_4a96edb8_(bus_4a96edb8_));
resized_LH1_xy_stateVar_Out1MaxTokenIndex resized_LH1_xy_stateVar_Out1MaxTokenIndex_1(.bus_344cf808_(CLK), 
  .bus_2e472a30_(bus_67d19bcd_), .bus_463825f8_(scheduler_u271), .bus_02e6a7a9_(scheduler_u272), 
  .bus_7668b64d_(bus_7668b64d_));
resized_LH1_xy_stateVar_rowRepeated resized_LH1_xy_stateVar_rowRepeated_1(.bus_1d013d35_(CLK), 
  .bus_1beb5227_(bus_67d19bcd_), .bus_0469fc4f_(repeatRowExpanded), .bus_51ae933d_(repeatRowExpanded_u24), 
  .bus_6a8dff02_(reset), .bus_733d2b23_(16'h1), .bus_70ada90a_(bus_70ada90a_));
resized_LH1_xy_structuralmemory_6d20861d_ resized_LH1_xy_structuralmemory_6d20861d__1(.CLK_u18(CLK), 
  .bus_28d40cb2_(bus_67d19bcd_), .bus_53538a8e_(bus_1c368516_), .bus_670f04d2_(3'h1), 
  .bus_5f174387_(bus_44b70675_), .bus_3aeafa89_(bus_178082e9_), .bus_10b1614e_(bus_17060ee9_), 
  .bus_2d676b21_(bus_2d676b21_), .bus_6bc2d2f4_(bus_6bc2d2f4_));
resized_LH1_xy_consumeRow resized_LH1_xy_consumeRow_instance(.CLK(CLK), .RESET(bus_67d19bcd_), 
  .GO(consumeRow_go), .port_6e9d7dff_(bus_72d7955d_), .port_33a398fc_(bus_7232d2ee_), 
  .port_2b507d31_(bus_1823b71b_), .port_58d4b229_(In1_DATA), .DONE(resized_LH1_xy_consumeRow_instance_DONE), 
  .RESULT(consumeRow), .RESULT_u1881(consumeRow_u30), .RESULT_u1886(consumeRow_u31), 
  .RESULT_u1887(consumeRow_u32), .RESULT_u1888(consumeRow_u33), .RESULT_u1889(consumeRow_u34), 
  .RESULT_u1882(consumeRow_u35), .RESULT_u1883(consumeRow_u36), .RESULT_u1884(consumeRow_u37), 
  .RESULT_u1885(consumeRow_u38), .RESULT_u1890(consumeRow_u39));
endmodule



module resized_LH1_xy_Kicker_43(CLK, RESET, bus_146eb89f_);
input		CLK;
input		RESET;
output		bus_146eb89f_;
reg		kicker_2=1'h0;
wire		bus_70d3cc08_;
wire		bus_16d87a23_;
reg		kicker_res=1'h0;
reg		kicker_1=1'h0;
wire		bus_7e1e6849_;
wire		bus_17e4289c_;
always @(posedge CLK)
begin
kicker_2<=bus_16d87a23_;
end
assign bus_70d3cc08_=~RESET;
assign bus_16d87a23_=bus_70d3cc08_&kicker_1;
always @(posedge CLK)
begin
kicker_res<=bus_17e4289c_;
end
always @(posedge CLK)
begin
kicker_1<=bus_70d3cc08_;
end
assign bus_7e1e6849_=~kicker_2;
assign bus_146eb89f_=kicker_res;
assign bus_17e4289c_=kicker_1&bus_70d3cc08_&bus_7e1e6849_;
endmodule



module resized_LH1_xy_forge_memory_512x16_33(CLK, EN, WE, ADDR, DIN, DOUT, DONE);
input		CLK;
input		EN;
input		WE;
input	[31:0]	ADDR;
input	[15:0]	DIN;
output	[15:0]	DOUT;
output		DONE;
wire		we_0;
wire	[15:0]	pre_dout_0;
wire		we_1;
wire	[15:0]	pre_dout_1;
wire		we_2;
wire	[15:0]	pre_dout_2;
wire		we_3;
wire	[15:0]	pre_dout_3;
reg	[15:0]	mux_out;
reg		wen_done;
assign we_0=WE&(ADDR[31:7]==25'h0);
assign we_1=WE&(ADDR[31:7]==25'h1);
assign we_2=WE&(ADDR[31:7]==25'h2);
assign we_3=WE&(ADDR[31:7]==25'h3);
always @(ADDR or pre_dout_0 or pre_dout_1 or pre_dout_2 or pre_dout_3)
begin
case (ADDR[31:7])25'd0:mux_out=pre_dout_0;
25'd1:mux_out=pre_dout_1;
25'd2:mux_out=pre_dout_2;
25'd3:mux_out=pre_dout_3;
default:mux_out=16'h0;
endcase end
always @(posedge CLK)
begin
wen_done<=WE;
end
assign DOUT=mux_out;
assign DONE=EN&!WE|wen_done;
//  Memory array element: COL: 0, ROW: 0
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_192(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[0]), .O(pre_dout_0[0]));
//  Memory array element: COL: 0, ROW: 1
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_193(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[1]), .O(pre_dout_0[1]));
//  Memory array element: COL: 0, ROW: 2
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_194(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[2]), .O(pre_dout_0[2]));
//  Memory array element: COL: 0, ROW: 3
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_195(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[3]), .O(pre_dout_0[3]));
//  Memory array element: COL: 0, ROW: 4
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_196(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[4]), .O(pre_dout_0[4]));
//  Memory array element: COL: 0, ROW: 5
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_197(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[5]), .O(pre_dout_0[5]));
//  Memory array element: COL: 0, ROW: 6
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_198(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[6]), .O(pre_dout_0[6]));
//  Memory array element: COL: 0, ROW: 7
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_199(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[7]), .O(pre_dout_0[7]));
//  Memory array element: COL: 0, ROW: 8
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_200(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[8]), .O(pre_dout_0[8]));
//  Memory array element: COL: 0, ROW: 9
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_201(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[9]), .O(pre_dout_0[9]));
//  Memory array element: COL: 0, ROW: 10
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_202(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[10]), .O(pre_dout_0[10]));
//  Memory array element: COL: 0, ROW: 11
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_203(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[11]), .O(pre_dout_0[11]));
//  Memory array element: COL: 0, ROW: 12
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_204(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[12]), .O(pre_dout_0[12]));
//  Memory array element: COL: 0, ROW: 13
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_205(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[13]), .O(pre_dout_0[13]));
//  Memory array element: COL: 0, ROW: 14
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_206(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[14]), .O(pre_dout_0[14]));
//  Memory array element: COL: 0, ROW: 15
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_207(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[15]), .O(pre_dout_0[15]));
//  Memory array element: COL: 1, ROW: 0
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_208(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[0]), .O(pre_dout_1[0]));
//  Memory array element: COL: 1, ROW: 1
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_209(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[1]), .O(pre_dout_1[1]));
//  Memory array element: COL: 1, ROW: 2
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_210(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[2]), .O(pre_dout_1[2]));
//  Memory array element: COL: 1, ROW: 3
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_211(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[3]), .O(pre_dout_1[3]));
//  Memory array element: COL: 1, ROW: 4
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_212(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[4]), .O(pre_dout_1[4]));
//  Memory array element: COL: 1, ROW: 5
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_213(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[5]), .O(pre_dout_1[5]));
//  Memory array element: COL: 1, ROW: 6
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_214(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[6]), .O(pre_dout_1[6]));
//  Memory array element: COL: 1, ROW: 7
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_215(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[7]), .O(pre_dout_1[7]));
//  Memory array element: COL: 1, ROW: 8
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_216(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[8]), .O(pre_dout_1[8]));
//  Memory array element: COL: 1, ROW: 9
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_217(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[9]), .O(pre_dout_1[9]));
//  Memory array element: COL: 1, ROW: 10
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_218(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[10]), .O(pre_dout_1[10]));
//  Memory array element: COL: 1, ROW: 11
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_219(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[11]), .O(pre_dout_1[11]));
//  Memory array element: COL: 1, ROW: 12
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_220(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[12]), .O(pre_dout_1[12]));
//  Memory array element: COL: 1, ROW: 13
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_221(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[13]), .O(pre_dout_1[13]));
//  Memory array element: COL: 1, ROW: 14
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_222(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[14]), .O(pre_dout_1[14]));
//  Memory array element: COL: 1, ROW: 15
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_223(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[15]), .O(pre_dout_1[15]));
//  Memory array element: COL: 2, ROW: 0
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_224(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[0]), .O(pre_dout_2[0]));
//  Memory array element: COL: 2, ROW: 1
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_225(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[1]), .O(pre_dout_2[1]));
//  Memory array element: COL: 2, ROW: 2
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_226(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[2]), .O(pre_dout_2[2]));
//  Memory array element: COL: 2, ROW: 3
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_227(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[3]), .O(pre_dout_2[3]));
//  Memory array element: COL: 2, ROW: 4
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_228(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[4]), .O(pre_dout_2[4]));
//  Memory array element: COL: 2, ROW: 5
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_229(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[5]), .O(pre_dout_2[5]));
//  Memory array element: COL: 2, ROW: 6
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_230(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[6]), .O(pre_dout_2[6]));
//  Memory array element: COL: 2, ROW: 7
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_231(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[7]), .O(pre_dout_2[7]));
//  Memory array element: COL: 2, ROW: 8
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_232(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[8]), .O(pre_dout_2[8]));
//  Memory array element: COL: 2, ROW: 9
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_233(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[9]), .O(pre_dout_2[9]));
//  Memory array element: COL: 2, ROW: 10
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_234(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[10]), .O(pre_dout_2[10]));
//  Memory array element: COL: 2, ROW: 11
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_235(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[11]), .O(pre_dout_2[11]));
//  Memory array element: COL: 2, ROW: 12
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_236(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[12]), .O(pre_dout_2[12]));
//  Memory array element: COL: 2, ROW: 13
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_237(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[13]), .O(pre_dout_2[13]));
//  Memory array element: COL: 2, ROW: 14
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_238(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[14]), .O(pre_dout_2[14]));
//  Memory array element: COL: 2, ROW: 15
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_239(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[15]), .O(pre_dout_2[15]));
//  Memory array element: COL: 3, ROW: 0
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_240(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[0]), .O(pre_dout_3[0]));
//  Memory array element: COL: 3, ROW: 1
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_241(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[1]), .O(pre_dout_3[1]));
//  Memory array element: COL: 3, ROW: 2
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_242(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[2]), .O(pre_dout_3[2]));
//  Memory array element: COL: 3, ROW: 3
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_243(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[3]), .O(pre_dout_3[3]));
//  Memory array element: COL: 3, ROW: 4
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_244(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[4]), .O(pre_dout_3[4]));
//  Memory array element: COL: 3, ROW: 5
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_245(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[5]), .O(pre_dout_3[5]));
//  Memory array element: COL: 3, ROW: 6
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_246(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[6]), .O(pre_dout_3[6]));
//  Memory array element: COL: 3, ROW: 7
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_247(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[7]), .O(pre_dout_3[7]));
//  Memory array element: COL: 3, ROW: 8
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_248(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[8]), .O(pre_dout_3[8]));
//  Memory array element: COL: 3, ROW: 9
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_249(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[9]), .O(pre_dout_3[9]));
//  Memory array element: COL: 3, ROW: 10
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_250(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[10]), .O(pre_dout_3[10]));
//  Memory array element: COL: 3, ROW: 11
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_251(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[11]), .O(pre_dout_3[11]));
//  Memory array element: COL: 3, ROW: 12
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_252(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[12]), .O(pre_dout_3[12]));
//  Memory array element: COL: 3, ROW: 13
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_253(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[13]), .O(pre_dout_3[13]));
//  Memory array element: COL: 3, ROW: 14
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_254(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[14]), .O(pre_dout_3[14]));
//  Memory array element: COL: 3, ROW: 15
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_255(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[15]), .O(pre_dout_3[15]));
endmodule



module resized_LH1_xy_structuralmemory_2108298e_(CLK_u17, bus_3a8ce0e8_, bus_32b68420_, bus_4efd6486_, bus_677fabb8_, bus_1c42c4da_, bus_5d26b9a7_, bus_37dd7726_, bus_0fe08b68_);
input		CLK_u17;
input		bus_3a8ce0e8_;
input	[31:0]	bus_32b68420_;
input	[2:0]	bus_4efd6486_;
input		bus_677fabb8_;
input		bus_1c42c4da_;
input	[15:0]	bus_5d26b9a7_;
output	[15:0]	bus_37dd7726_;
output		bus_0fe08b68_;
wire		not_6d5e0bde_u0;
wire		or_696ea22a_u0;
wire		or_0a807e88_u0;
wire	[15:0]	bus_3af7f7e9_;
wire		and_1724ad36_u0;
reg		logicalMem_9baf256_we_delay0_u0=1'h0;
assign not_6d5e0bde_u0=~bus_1c42c4da_;
assign or_696ea22a_u0=bus_677fabb8_|bus_1c42c4da_;
assign or_0a807e88_u0=and_1724ad36_u0|logicalMem_9baf256_we_delay0_u0;
resized_LH1_xy_forge_memory_512x16_33 resized_LH1_xy_forge_memory_512x16_33_instance0(.CLK(CLK_u17), 
  .EN(or_696ea22a_u0), .WE(bus_1c42c4da_), .ADDR(bus_32b68420_), .DIN(bus_5d26b9a7_), 
  .DOUT(bus_3af7f7e9_), .DONE());
assign and_1724ad36_u0=bus_677fabb8_&not_6d5e0bde_u0;
always @(posedge CLK_u17 or posedge bus_3a8ce0e8_)
begin
if (bus_3a8ce0e8_)
logicalMem_9baf256_we_delay0_u0<=1'h0;
else logicalMem_9baf256_we_delay0_u0<=bus_1c42c4da_;
end
assign bus_37dd7726_=bus_3af7f7e9_;
assign bus_0fe08b68_=or_0a807e88_u0;
endmodule



module resized_LH1_xy_stateVar_Out1PortEnable(bus_7dadb443_, bus_2cfd1fd9_, bus_105e9f86_, bus_4406fa74_, bus_2698717b_);
input		bus_7dadb443_;
input		bus_2cfd1fd9_;
input		bus_105e9f86_;
input		bus_4406fa74_;
output		bus_2698717b_;
reg		stateVar_Out1PortEnable_u3=1'h0;
assign bus_2698717b_=stateVar_Out1PortEnable_u3;
always @(posedge bus_7dadb443_ or posedge bus_2cfd1fd9_)
begin
if (bus_2cfd1fd9_)
stateVar_Out1PortEnable_u3<=1'h0;
else if (bus_105e9f86_)
stateVar_Out1PortEnable_u3<=bus_4406fa74_;
end
endmodule



module resized_LH1_xy_endianswapper_294583ce_(endianswapper_294583ce_in, endianswapper_294583ce_out);
input	[15:0]	endianswapper_294583ce_in;
output	[15:0]	endianswapper_294583ce_out;
assign endianswapper_294583ce_out=endianswapper_294583ce_in;
endmodule



module resized_LH1_xy_endianswapper_449ee5a2_(endianswapper_449ee5a2_in, endianswapper_449ee5a2_out);
input	[15:0]	endianswapper_449ee5a2_in;
output	[15:0]	endianswapper_449ee5a2_out;
assign endianswapper_449ee5a2_out=endianswapper_449ee5a2_in;
endmodule



module resized_LH1_xy_stateVar_x(bus_78bae313_, bus_6b0a580d_, bus_4a98ed23_, bus_5ce6cb87_, bus_3e718195_, bus_18105192_, bus_72d7955d_);
input		bus_78bae313_;
input		bus_6b0a580d_;
input		bus_4a98ed23_;
input	[15:0]	bus_5ce6cb87_;
input		bus_3e718195_;
input	[15:0]	bus_18105192_;
output	[15:0]	bus_72d7955d_;
reg	[15:0]	stateVar_x_u3=16'h0;
wire	[15:0]	mux_30d4a5a6_u0;
wire		or_3b129db7_u0;
wire	[15:0]	endianswapper_294583ce_out;
wire	[15:0]	endianswapper_449ee5a2_out;
always @(posedge bus_78bae313_ or posedge bus_6b0a580d_)
begin
if (bus_6b0a580d_)
stateVar_x_u3<=16'h0;
else if (or_3b129db7_u0)
stateVar_x_u3<=endianswapper_449ee5a2_out;
end
assign mux_30d4a5a6_u0=(bus_4a98ed23_)?bus_5ce6cb87_:16'h0;
assign or_3b129db7_u0=bus_4a98ed23_|bus_3e718195_;
resized_LH1_xy_endianswapper_294583ce_ resized_LH1_xy_endianswapper_294583ce__1(.endianswapper_294583ce_in(stateVar_x_u3), 
  .endianswapper_294583ce_out(endianswapper_294583ce_out));
resized_LH1_xy_endianswapper_449ee5a2_ resized_LH1_xy_endianswapper_449ee5a2__1(.endianswapper_449ee5a2_in(mux_30d4a5a6_u0), 
  .endianswapper_449ee5a2_out(endianswapper_449ee5a2_out));
assign bus_72d7955d_=endianswapper_294583ce_out;
endmodule



module resized_LH1_xy_globalreset_physical_790ef242_(bus_664d27ed_, bus_42d18000_, bus_67d19bcd_);
input		bus_664d27ed_;
input		bus_42d18000_;
output		bus_67d19bcd_;
wire		not_335af6fb_u0;
wire		or_3e6c814d_u0;
wire		and_38eec71d_u0;
reg		sample_u39=1'h0;
reg		cross_u39=1'h0;
reg		final_u39=1'h1;
reg		glitch_u39=1'h0;
assign not_335af6fb_u0=~and_38eec71d_u0;
assign or_3e6c814d_u0=bus_42d18000_|final_u39;
assign and_38eec71d_u0=cross_u39&glitch_u39;
always @(posedge bus_664d27ed_)
begin
sample_u39<=1'h1;
end
always @(posedge bus_664d27ed_)
begin
cross_u39<=sample_u39;
end
assign bus_67d19bcd_=or_3e6c814d_u0;
always @(posedge bus_664d27ed_)
begin
final_u39<=not_335af6fb_u0;
end
always @(posedge bus_664d27ed_)
begin
glitch_u39<=cross_u39;
end
endmodule



module resized_LH1_xy_endianswapper_50e686b7_(endianswapper_50e686b7_in, endianswapper_50e686b7_out);
input	[31:0]	endianswapper_50e686b7_in;
output	[31:0]	endianswapper_50e686b7_out;
assign endianswapper_50e686b7_out=32'h0;
endmodule



module resized_LH1_xy_endianswapper_5eaf9e01_(endianswapper_5eaf9e01_in, endianswapper_5eaf9e01_out);
input	[31:0]	endianswapper_5eaf9e01_in;
output	[31:0]	endianswapper_5eaf9e01_out;
assign endianswapper_5eaf9e01_out=32'h0;
endmodule



module resized_LH1_xy_stateVar_fsmOldState_resized_LH1_xy(bus_201216da_, bus_66f3f92d_, bus_7673123e_, bus_3fa4cd9c_, bus_3d2b1c2b_);
input		bus_201216da_;
input		bus_66f3f92d_;
input		bus_7673123e_;
input	[31:0]	bus_3fa4cd9c_;
output	[31:0]	bus_3d2b1c2b_;
wire	[31:0]	endianswapper_50e686b7_out;
wire	[31:0]	endianswapper_5eaf9e01_out;
resized_LH1_xy_endianswapper_50e686b7_ resized_LH1_xy_endianswapper_50e686b7__1(.endianswapper_50e686b7_in(32'h0), 
  .endianswapper_50e686b7_out(endianswapper_50e686b7_out));
assign bus_3d2b1c2b_=32'h0;
resized_LH1_xy_endianswapper_5eaf9e01_ resized_LH1_xy_endianswapper_5eaf9e01__1(.endianswapper_5eaf9e01_in(32'h0), 
  .endianswapper_5eaf9e01_out(endianswapper_5eaf9e01_out));
endmodule



module resized_LH1_xy_reset(CLK, RESET, GO, RESULT, RESULT_u1852, RESULT_u1853, RESULT_u1854, DONE);
input		CLK;
input		RESET;
input		GO;
output		RESULT;
output	[15:0]	RESULT_u1852;
output		RESULT_u1853;
output	[15:0]	RESULT_u1854;
output		DONE;
reg		reg_3ad0296b_u0=1'h0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3ad0296b_u0<=1'h0;
else reg_3ad0296b_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u1852=16'h1;
assign RESULT_u1853=GO;
assign RESULT_u1854=16'h0;
assign DONE=reg_3ad0296b_u0;
endmodule



module resized_LH1_xy_simplememoryreferee_07b85719_(bus_0b291028_, bus_154448d0_, bus_2afbec8d_, bus_1f157a32_, bus_6d609752_, bus_5486e989_, bus_25b9b8db_, bus_0756d9ea_, bus_588863ee_, bus_79191f33_, bus_4bdb631c_, bus_043f5796_, bus_0dea0337_, bus_47674f00_, bus_41a72575_, bus_54d5acc6_, bus_1823b71b_, bus_5d969c8b_, bus_053c348c_);
input		bus_0b291028_;
input		bus_154448d0_;
input		bus_2afbec8d_;
input	[15:0]	bus_1f157a32_;
input		bus_6d609752_;
input	[15:0]	bus_5486e989_;
input	[31:0]	bus_25b9b8db_;
input	[2:0]	bus_0756d9ea_;
input		bus_588863ee_;
input	[31:0]	bus_79191f33_;
input	[2:0]	bus_4bdb631c_;
output	[15:0]	bus_043f5796_;
output	[31:0]	bus_0dea0337_;
output		bus_47674f00_;
output		bus_41a72575_;
output	[2:0]	bus_54d5acc6_;
output		bus_1823b71b_;
output	[15:0]	bus_5d969c8b_;
output		bus_053c348c_;
wire		and_3da3be87_u0;
wire		not_6d00abe4_u0;
wire	[15:0]	mux_31582b13_u0;
reg		done_qual_u165=1'h0;
reg		done_qual_u166_u0=1'h0;
wire		or_2ce40357_u0;
wire		or_6c4eb6fa_u0;
wire		and_004ab45d_u0;
wire		or_343d2925_u0;
wire		not_0bcfe976_u0;
wire	[31:0]	mux_1ee5a43a_u0;
assign and_3da3be87_u0=or_2ce40357_u0&bus_2afbec8d_;
assign not_6d00abe4_u0=~bus_2afbec8d_;
assign mux_31582b13_u0=({16{bus_6d609752_}}&bus_5486e989_);
always @(posedge bus_0b291028_)
begin
if (bus_154448d0_)
done_qual_u165<=1'h0;
else done_qual_u165<=bus_6d609752_;
end
always @(posedge bus_0b291028_)
begin
if (bus_154448d0_)
done_qual_u166_u0<=1'h0;
else done_qual_u166_u0<=bus_588863ee_;
end
assign or_2ce40357_u0=bus_588863ee_|done_qual_u166_u0;
assign or_6c4eb6fa_u0=bus_6d609752_|done_qual_u165;
assign and_004ab45d_u0=or_6c4eb6fa_u0&bus_2afbec8d_;
assign or_343d2925_u0=bus_6d609752_|bus_588863ee_;
assign not_0bcfe976_u0=~bus_2afbec8d_;
assign bus_043f5796_=mux_31582b13_u0;
assign bus_0dea0337_=mux_1ee5a43a_u0;
assign bus_47674f00_=bus_6d609752_;
assign bus_41a72575_=or_343d2925_u0;
assign bus_54d5acc6_=3'h1;
assign bus_1823b71b_=and_004ab45d_u0;
assign bus_5d969c8b_=bus_1f157a32_;
assign bus_053c348c_=and_3da3be87_u0;
assign mux_1ee5a43a_u0=(bus_6d609752_)?bus_25b9b8db_:bus_79191f33_;
endmodule



module resized_LH1_xy_endianswapper_1917bc44_(endianswapper_1917bc44_in, endianswapper_1917bc44_out);
input		endianswapper_1917bc44_in;
output		endianswapper_1917bc44_out;
assign endianswapper_1917bc44_out=endianswapper_1917bc44_in;
endmodule



module resized_LH1_xy_endianswapper_52feac5d_(endianswapper_52feac5d_in, endianswapper_52feac5d_out);
input		endianswapper_52feac5d_in;
output		endianswapper_52feac5d_out;
assign endianswapper_52feac5d_out=endianswapper_52feac5d_in;
endmodule



module resized_LH1_xy_stateVar_fsmState_resized_LH1_xy(bus_3631bc0b_, bus_0708d8fb_, bus_4602c2a7_, bus_3c662fde_, bus_382ad4dd_);
input		bus_3631bc0b_;
input		bus_0708d8fb_;
input		bus_4602c2a7_;
input		bus_3c662fde_;
output		bus_382ad4dd_;
wire		endianswapper_1917bc44_out;
wire		endianswapper_52feac5d_out;
reg		stateVar_fsmState_resized_LH1_xy_u0=1'h0;
resized_LH1_xy_endianswapper_1917bc44_ resized_LH1_xy_endianswapper_1917bc44__1(.endianswapper_1917bc44_in(bus_3c662fde_), 
  .endianswapper_1917bc44_out(endianswapper_1917bc44_out));
resized_LH1_xy_endianswapper_52feac5d_ resized_LH1_xy_endianswapper_52feac5d__1(.endianswapper_52feac5d_in(stateVar_fsmState_resized_LH1_xy_u0), 
  .endianswapper_52feac5d_out(endianswapper_52feac5d_out));
assign bus_382ad4dd_=endianswapper_52feac5d_out;
always @(posedge bus_3631bc0b_ or posedge bus_0708d8fb_)
begin
if (bus_0708d8fb_)
stateVar_fsmState_resized_LH1_xy_u0<=1'h0;
else if (bus_4602c2a7_)
stateVar_fsmState_resized_LH1_xy_u0<=endianswapper_1917bc44_out;
end
endmodule



module resized_LH1_xy_repeatRowExpanded(CLK, RESET, GO, port_1819de90_, port_5d43c181_, port_00ba0d3b_, port_6635e8af_, RESULT, RESULT_u1855, RESULT_u1856, RESULT_u1857, RESULT_u1858, RESULT_u1859, RESULT_u1860, RESULT_u1861, RESULT_u1862, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_1819de90_;
input		port_5d43c181_;
input	[15:0]	port_00ba0d3b_;
input		port_6635e8af_;
output		RESULT;
output	[15:0]	RESULT_u1855;
output		RESULT_u1856;
output	[31:0]	RESULT_u1857;
output	[2:0]	RESULT_u1858;
output		RESULT_u1859;
output	[31:0]	RESULT_u1860;
output	[15:0]	RESULT_u1861;
output	[2:0]	RESULT_u1862;
output		DONE;
wire	[15:0]	add;
wire		and_u3134_u0;
wire signed	[31:0]	lessThan_a_signed;
wire signed	[31:0]	lessThan_b_signed;
wire		lessThan;
wire		and_u3135_u0;
wire		and_u3136_u0;
wire		not_u525_u0;
reg		and_delayed_u206=1'h0;
wire	[31:0]	add_u371;
wire		and_u3137_u0;
wire	[31:0]	add_u372;
reg		reg_5b526fb2_u0=1'h0;
wire		and_u3138_u0;
wire		or_u893_u0;
wire	[31:0]	add_u373;
reg	[31:0]	syncEnable_u549=32'h0;
wire		and_u3139_u0;
wire	[31:0]	mux_u314;
wire		or_u894_u0;
reg		reg_02223f9e_u0=1'h0;
assign add=port_1819de90_+16'h1;
assign and_u3134_u0=and_u3135_u0&or_u894_u0;
assign lessThan_a_signed=mux_u314;
assign lessThan_b_signed=32'h200;
assign lessThan=lessThan_a_signed<lessThan_b_signed;
assign and_u3135_u0=or_u894_u0&lessThan;
assign and_u3136_u0=or_u894_u0&not_u525_u0;
assign not_u525_u0=~lessThan;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u206<=1'h0;
else and_delayed_u206<=and_u3134_u0;
end
assign add_u371=mux_u314+32'h0;
assign and_u3137_u0=and_u3134_u0&port_5d43c181_;
assign add_u372=mux_u314+32'h0;
always @(posedge CLK or posedge and_u3134_u0 or posedge or_u893_u0)
begin
if (or_u893_u0)
reg_5b526fb2_u0<=1'h0;
else if (and_u3134_u0)
reg_5b526fb2_u0<=1'h1;
else reg_5b526fb2_u0<=reg_5b526fb2_u0;
end
assign and_u3138_u0=reg_5b526fb2_u0&port_6635e8af_;
assign or_u893_u0=and_u3138_u0|RESET;
assign add_u373=mux_u314+32'h1;
always @(posedge CLK)
begin
if (and_u3134_u0)
syncEnable_u549<=add_u373;
end
assign and_u3139_u0=and_u3136_u0&or_u894_u0;
assign mux_u314=(reg_02223f9e_u0)?32'h0:syncEnable_u549;
assign or_u894_u0=reg_02223f9e_u0|and_delayed_u206;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_02223f9e_u0<=1'h0;
else reg_02223f9e_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u1855=add;
assign RESULT_u1856=and_u3134_u0;
assign RESULT_u1857=add_u371;
assign RESULT_u1858=3'h1;
assign RESULT_u1859=and_u3134_u0;
assign RESULT_u1860=add_u372;
assign RESULT_u1861=port_00ba0d3b_;
assign RESULT_u1862=3'h1;
assign DONE=and_u3139_u0;
endmodule



module resized_LH1_xy_simplememoryreferee_4f8eca27_(bus_13a35abe_, bus_537d7f21_, bus_67df8591_, bus_26c151a5_, bus_7e206820_, bus_0bdb3367_, bus_3ac51013_, bus_7de908f2_, bus_2043bfd1_, bus_0ca641af_, bus_6077dae8_, bus_0fd5a0d9_, bus_2444a5e9_, bus_242bf648_, bus_528d16c5_, bus_17060ee9_, bus_1c368516_, bus_178082e9_, bus_44b70675_, bus_527ad470_, bus_7232d2ee_, bus_6818c058_, bus_0af0ab39_, bus_7cc52ea4_);
input		bus_13a35abe_;
input		bus_537d7f21_;
input		bus_67df8591_;
input	[15:0]	bus_26c151a5_;
input		bus_7e206820_;
input	[15:0]	bus_0bdb3367_;
input	[31:0]	bus_3ac51013_;
input	[2:0]	bus_7de908f2_;
input		bus_2043bfd1_;
input	[15:0]	bus_0ca641af_;
input	[31:0]	bus_6077dae8_;
input	[2:0]	bus_0fd5a0d9_;
input		bus_2444a5e9_;
input	[31:0]	bus_242bf648_;
input	[2:0]	bus_528d16c5_;
output	[15:0]	bus_17060ee9_;
output	[31:0]	bus_1c368516_;
output		bus_178082e9_;
output		bus_44b70675_;
output	[2:0]	bus_527ad470_;
output		bus_7232d2ee_;
output		bus_6818c058_;
output	[15:0]	bus_0af0ab39_;
output		bus_7cc52ea4_;
wire		or_2f55f270_u0;
wire	[31:0]	mux_67b2c4f4_u0;
wire		or_41538c38_u0;
reg		done_qual_u167_u0=1'h0;
wire		not_64863029_u0;
wire		or_5e1e23ef_u0;
reg		done_qual_u168_u0=1'h0;
wire		not_0cda1e68_u0;
wire		and_2f0cb179_u0;
wire		and_4fbc91a9_u0;
wire		or_45dae622_u0;
reg		done_qual_u169_u0=1'h0;
wire		or_5851fc8c_u0;
wire	[15:0]	mux_452c4731_u0;
wire		and_6b9f5982_u0;
wire		not_120a84b4_u0;
assign or_2f55f270_u0=bus_7e206820_|done_qual_u168_u0;
assign mux_67b2c4f4_u0=({32{bus_7e206820_}}&bus_3ac51013_)|({32{bus_2043bfd1_}}&bus_6077dae8_)|({32{bus_2444a5e9_}}&bus_242bf648_);
assign or_41538c38_u0=bus_2444a5e9_|done_qual_u167_u0;
assign bus_17060ee9_=mux_452c4731_u0;
assign bus_1c368516_=mux_67b2c4f4_u0;
assign bus_178082e9_=or_5851fc8c_u0;
assign bus_44b70675_=or_5e1e23ef_u0;
assign bus_527ad470_=3'h1;
assign bus_7232d2ee_=and_6b9f5982_u0;
assign bus_6818c058_=and_2f0cb179_u0;
assign bus_0af0ab39_=bus_26c151a5_;
assign bus_7cc52ea4_=and_4fbc91a9_u0;
always @(posedge bus_13a35abe_)
begin
if (bus_537d7f21_)
done_qual_u167_u0<=1'h0;
else done_qual_u167_u0<=bus_2444a5e9_;
end
assign not_64863029_u0=~bus_67df8591_;
assign or_5e1e23ef_u0=bus_7e206820_|bus_2043bfd1_|bus_2444a5e9_;
always @(posedge bus_13a35abe_)
begin
if (bus_537d7f21_)
done_qual_u168_u0<=1'h0;
else done_qual_u168_u0<=bus_7e206820_;
end
assign not_0cda1e68_u0=~bus_67df8591_;
assign and_2f0cb179_u0=or_45dae622_u0&bus_67df8591_;
assign and_4fbc91a9_u0=or_41538c38_u0&bus_67df8591_;
assign or_45dae622_u0=bus_2043bfd1_|done_qual_u169_u0;
always @(posedge bus_13a35abe_)
begin
if (bus_537d7f21_)
done_qual_u169_u0<=1'h0;
else done_qual_u169_u0<=bus_2043bfd1_;
end
assign or_5851fc8c_u0=bus_7e206820_|bus_2043bfd1_;
assign mux_452c4731_u0=(bus_7e206820_)?bus_0bdb3367_:bus_0ca641af_;
assign and_6b9f5982_u0=or_2f55f270_u0&bus_67df8591_;
assign not_120a84b4_u0=~bus_67df8591_;
endmodule



module resized_LH1_xy_scheduler(CLK, RESET, GO, port_6105e58c_, port_0a81f2c6_, port_3bb784d0_, port_1ca215c6_, port_5071c1a7_, port_008a440f_, port_1ba874b3_, port_63d562ec_, port_2ccab656_, port_2adbeb14_, port_218764d5_, port_51b44ade_, port_58303e5a_, port_1be35c61_, RESULT, RESULT_u1863, RESULT_u1864, RESULT_u1865, RESULT_u1866, RESULT_u1867, RESULT_u1868, RESULT_u1869, RESULT_u1870, RESULT_u1871, RESULT_u1872, RESULT_u1873, RESULT_u1874, RESULT_u1875, RESULT_u1876, RESULT_u1877, RESULT_u1878, RESULT_u1879, RESULT_u1880, DONE);
input		CLK;
input		RESET;
input		GO;
input	[31:0]	port_6105e58c_;
input		port_0a81f2c6_;
input	[31:0]	port_3bb784d0_;
input	[31:0]	port_1ca215c6_;
input		port_5071c1a7_;
input	[15:0]	port_008a440f_;
input	[15:0]	port_1ba874b3_;
input		port_63d562ec_;
input	[15:0]	port_2ccab656_;
input		port_2adbeb14_;
input		port_218764d5_;
input		port_51b44ade_;
input		port_58303e5a_;
input		port_1be35c61_;
output		RESULT;
output	[31:0]	RESULT_u1863;
output		RESULT_u1864;
output		RESULT_u1865;
output		RESULT_u1866;
output	[31:0]	RESULT_u1867;
output		RESULT_u1868;
output	[31:0]	RESULT_u1869;
output		RESULT_u1870;
output		RESULT_u1871;
output		RESULT_u1872;
output	[31:0]	RESULT_u1873;
output	[2:0]	RESULT_u1874;
output		RESULT_u1875;
output	[15:0]	RESULT_u1876;
output		RESULT_u1877;
output		RESULT_u1878;
output	[15:0]	RESULT_u1879;
output		RESULT_u1880;
output		DONE;
wire		and_u3140_u0;
wire		lessThan;
wire	[15:0]	lessThan_b_unsigned;
wire	[15:0]	lessThan_a_unsigned;
wire	[15:0]	equals_a_unsigned;
wire	[15:0]	equals_b_unsigned;
wire		equals;
wire	[15:0]	lessThan_u74_a_unsigned;
wire		lessThan_u74;
wire	[15:0]	lessThan_u74_b_unsigned;
wire		andOp;
wire	[15:0]	equals_u164_a_unsigned;
wire		equals_u164;
wire	[15:0]	equals_u164_b_unsigned;
wire		equals_u165;
wire signed	[31:0]	equals_u165_a_signed;
wire signed	[31:0]	equals_u165_b_signed;
wire		not_u526_u0;
wire		and_u3141_u0;
wire		and_u3142_u0;
wire		andOp_u173;
wire		and_u3143_u0;
wire		and_u3144_u0;
wire		not_u527_u0;
wire		simplePinWrite;
wire		and_u3145_u0;
wire		not_u528_u0;
wire		and_u3146_u0;
wire		simplePinWrite_u466;
wire		and_u3147_u0;
wire		not_u529_u0;
wire		and_u3148_u0;
wire		simplePinWrite_u467;
wire		and_u3149_u0;
reg		reg_297a657a_u0=1'h0;
reg		reg_378e778c_u0=1'h0;
reg		reg_50917495_u0=1'h0;
reg		reg_05074d01_u0=1'h0;
reg		reg_2c3cec3a_u0=1'h0;
reg		reg_7bc1bfcd_u0=1'h0;
reg		reg_77047715_u0=1'h0;
reg		reg_6fbb03a9_u0=1'h0;
reg		reg_401b0405_u0=1'h0;
reg		reg_5b15db0b_u0=1'h0;
reg		reg_5c74f06b_u0=1'h0;
reg		reg_2ecaeed5_u0=1'h0;
reg		reg_64fa00de_u0=1'h0;
reg		reg_65acfd8b_u0=1'h0;
reg		reg_2cb89c91_u0=1'h0;
reg		reg_4e012e31_u0=1'h0;
reg		reg_324e3a7d_u0=1'h0;
reg		reg_324e3a7d_result_delayed_u0=1'h0;
reg		reg_1a7a9643_u0=1'h0;
reg		reg_40d160ea_u0=1'h0;
reg		reg_05c10dfa_u0=1'h0;
reg		reg_357b5d40_u0=1'h0;
reg		reg_1b8047bd_u0=1'h0;
reg		reg_6d5cb91c_u0=1'h0;
reg		reg_5f68d729_u0=1'h0;
reg		reg_2d3a4979_u0=1'h0;
reg		reg_258519cc_u0=1'h0;
reg		reg_7b23ef69_u0=1'h0;
reg		reg_4e9c06d0_u0=1'h0;
reg		reg_710c3541_u0=1'h0;
reg		reg_6e5ada14_u0=1'h0;
reg		reg_030c675e_u0=1'h0;
reg		reg_2139e56a_u0=1'h0;
reg		reg_01aa19f9_u0=1'h0;
reg		reg_00bce4e8_u0=1'h0;
reg		reg_1de599bc_u0=1'h0;
reg		reg_79b769ec_u0=1'h0;
reg		reg_17e75387_u0=1'h0;
reg		reg_689528f4_u0=1'h0;
reg		reg_3e784e1c_u0=1'h0;
reg		reg_387e0416_u0=1'h0;
reg		reg_43039f69_u0=1'h0;
reg		reg_6806d06c_u0=1'h0;
reg		reg_6b6d7306_u0=1'h0;
reg		reg_138117ea_u0=1'h0;
reg		reg_683a6054_u0=1'h0;
reg		reg_5aa7d6c8_u0=1'h0;
reg		reg_05286558_u0=1'h0;
reg		reg_55180568_u0=1'h0;
reg		reg_71bdf9cc_u0=1'h0;
reg		reg_79b769ec_result_delayed_u0=1'h0;
reg		reg_3d4ff93c_u0=1'h0;
reg		reg_1b57bf2f_u0=1'h0;
reg		reg_33167b6e_u0=1'h0;
reg		reg_4b39e741_u0=1'h0;
reg		reg_63daa7a1_u0=1'h0;
reg		reg_3b4c4b37_u0=1'h0;
reg		reg_5e96aee9_u0=1'h0;
reg		reg_47eb2b6a_u0=1'h0;
reg		reg_09c6d144_u0=1'h0;
reg		reg_7ff55f76_u0=1'h0;
reg		reg_3c8b940e_u0=1'h0;
reg		reg_4e70c2f7_u0=1'h0;
reg		reg_6e5ada14_result_delayed_u0=1'h0;
reg		reg_3e784e1c_result_delayed_u0=1'h0;
reg		reg_638aaf04_u0=1'h0;
reg		reg_2c075897_u0=1'h0;
reg		reg_0a611af4_u0=1'h0;
reg		reg_49dd354a_u0=1'h0;
reg		reg_3212b28a_u0=1'h0;
reg		reg_66095291_u0=1'h0;
reg		reg_40adac30_u0=1'h0;
reg		reg_33b11310_u0=1'h0;
reg		reg_27e96f4d_u0=1'h0;
reg		reg_0a0626a2_u0=1'h0;
reg		reg_0edfde7a_u0=1'h0;
reg		reg_54826c24_u0=1'h0;
reg		reg_43039f69_result_delayed_u0=1'h0;
reg		reg_5780a32a_u0=1'h0;
reg		reg_63c2bf6e_u0=1'h0;
reg		reg_1f49a7e5_u0=1'h0;
reg		reg_63314f9f_u0=1'h0;
reg		reg_281f24ad_u0=1'h0;
reg		reg_3212b28a_result_delayed_u0=1'h0;
reg		reg_3f347781_u0=1'h0;
reg		reg_05fa154c_u0=1'h0;
wire		and_u3150_u0;
reg		reg_2139e56a_result_delayed_u0=1'h0;
reg		reg_107844c4_u0=1'h0;
reg		reg_318c1131_u0=1'h0;
reg		reg_689528f4_result_delayed_u0=1'h0;
reg		reg_32fe623a_u0=1'h0;
reg		reg_69fad53c_u0=1'h0;
reg		reg_35da391c_u0=1'h0;
reg		reg_23499f80_u0=1'h0;
reg		reg_2f7313b9_u0=1'h0;
reg		reg_2ecaeed5_result_delayed_u0=1'h0;
reg		reg_107844c4_result_delayed_u0=1'h0;
reg		reg_0bfe7f33_u0=1'h0;
reg		reg_7a51229e_u0=1'h0;
reg		reg_33167b6e_result_delayed_u0=1'h0;
reg		reg_6e8b025a_u0=1'h0;
reg		reg_546fd8be_u0=1'h0;
reg		reg_7a88ee59_u0=1'h0;
reg		reg_0c3478e6_u0=1'h0;
reg		reg_1de599bc_result_delayed_u0=1'h0;
reg		reg_05074d01_result_delayed_u0=1'h0;
reg		reg_1dd4f50d_u0=1'h0;
reg		reg_49f0052b_u0=1'h0;
reg		reg_7217fecc_u0=1'h0;
reg		reg_7e56828a_u0=1'h0;
reg		reg_32a6867b_u0=1'h0;
reg		reg_6dc4bd1b_u0=1'h0;
reg		reg_23b56b6a_u0=1'h0;
reg		reg_0edfde7a_result_delayed_u0=1'h0;
reg		reg_5f095be9_u0=1'h0;
reg		reg_43d5e336_u0=1'h0;
reg		reg_64fa00de_result_delayed_u0=1'h0;
reg		reg_01db913f_u0=1'h0;
reg		reg_355135b7_u0=1'h0;
reg		reg_429ea278_u0=1'h0;
reg		reg_6109ede1_u0=1'h0;
reg		reg_049d2474_u0=1'h0;
reg		reg_279d2f74_u0=1'h0;
reg		reg_536a7781_u0=1'h0;
reg		reg_7c5e48af_u0=1'h0;
reg		reg_355135b7_result_delayed_u0=1'h0;
reg		reg_03e66f15_u0=1'h0;
reg		reg_0a6e669d_u0=1'h0;
reg		reg_29259ddf_u0=1'h0;
reg		reg_14fc4001_u0=1'h0;
reg		reg_7c7f1881_u0=1'h0;
reg		reg_5a95fe6b_u0=1'h0;
reg		reg_52d98a27_u0=1'h0;
reg		reg_640558fa_u0=1'h0;
reg		reg_05c10dfa_result_delayed_u0=1'h0;
reg		reg_7b23ef69_result_delayed_u0=1'h0;
reg		reg_10dd85da_u0=1'h0;
reg		reg_6685c38c_u0=1'h0;
reg		reg_00326d3c_u0=1'h0;
reg		reg_65acfd8b_result_delayed_u0=1'h0;
reg		reg_12289738_u0=1'h0;
reg		reg_05fa154c_result_delayed_u0=1'h0;
reg		reg_4a292b3c_u0=1'h0;
reg		reg_5011c507_u0=1'h0;
reg		reg_3c99258f_u0=1'h0;
reg		reg_792a283d_u0=1'h0;
reg		reg_6a06c71e_u0=1'h0;
reg		reg_0c3478e6_result_delayed_u0=1'h0;
reg		reg_47f4e6ec_u0=1'h0;
reg		reg_32e22ff9_u0=1'h0;
reg		reg_1ca67dbd_u0=1'h0;
reg		reg_3b393219_u0=1'h0;
reg		reg_0304da20_u0=1'h0;
reg		reg_40adac30_result_delayed_u0=1'h0;
reg		reg_6e43fb69_u0=1'h0;
reg		reg_5f7ee655_u0=1'h0;
reg		reg_0304da20_result_delayed_u0=1'h0;
reg		reg_60f891d5_u0=1'h0;
reg		reg_5eccd3e3_u0=1'h0;
reg		reg_04854db4_u0=1'h0;
reg		reg_6b6d7306_result_delayed_u0=1'h0;
reg		reg_41025437_u0=1'h0;
reg		reg_35ff7cc6_u0=1'h0;
reg		reg_437f3245_u0=1'h0;
reg		reg_1536c80b_u0=1'h0;
reg		reg_1536340b_u0=1'h0;
reg		reg_33167b6e_result_delayed_result_delayed_u0=1'h0;
reg		reg_6fc41285_u0=1'h0;
reg		reg_11d4a896_u0=1'h0;
reg		reg_32a6867b_result_delayed_u0=1'h0;
reg		reg_4e9c06d0_result_delayed_u0=1'h0;
reg		reg_1e58db1f_u0=1'h0;
reg		reg_74e3dda4_u0=1'h0;
reg		reg_7a3ed379_u0=1'h0;
reg		reg_2e62ff2a_u0=1'h0;
reg		reg_7a88ee59_result_delayed_u0=1'h0;
reg		reg_05074d01_result_delayed_result_delayed_u0=1'h0;
reg		reg_0319ee54_u0=1'h0;
reg		reg_4f8202d0_u0=1'h0;
reg		reg_2349ca1b_u0=1'h0;
reg		reg_7f7d622f_u0=1'h0;
reg		reg_6e8b025a_result_delayed_u0=1'h0;
reg		reg_2bfa4eac_u0=1'h0;
reg		reg_7e0ad75d_u0=1'h0;
reg		reg_7b23ef69_result_delayed_result_delayed_u0=1'h0;
reg		reg_1a836fd8_u0=1'h0;
reg		reg_342c7170_u0=1'h0;
reg		reg_69fad53c_result_delayed_u0=1'h0;
reg		reg_3622ef46_u0=1'h0;
reg		reg_261ccf7a_u0=1'h0;
reg		reg_6741a229_u0=1'h0;
reg		reg_29259ddf_result_delayed_u0=1'h0;
reg		reg_0fb3eac1_u0=1'h0;
reg		reg_75b844ca_u0=1'h0;
reg		reg_4d6a0c19_u0=1'h0;
reg		reg_281f24ad_result_delayed_u0=1'h0;
reg		reg_5c72dd07_u0=1'h0;
reg		reg_2c075897_result_delayed_u0=1'h0;
reg		reg_6c0ed978_u0=1'h0;
reg		reg_7106847e_u0=1'h0;
reg		reg_5cd43dad_u0=1'h0;
reg		reg_63ada2d0_u0=1'h0;
reg		reg_6812ad6d_u0=1'h0;
reg		reg_14fc4001_result_delayed_u0=1'h0;
reg		reg_3bc4d242_u0=1'h0;
reg		reg_47b1c63c_u0=1'h0;
reg		reg_2a1c2b8c_u0=1'h0;
reg		reg_1ab96b28_u0=1'h0;
reg		reg_60f891d5_result_delayed_u0=1'h0;
reg		reg_57713ae7_u0=1'h0;
reg		reg_2dbd2c2b_u0=1'h0;
reg		reg_682b29b0_u0=1'h0;
reg		reg_357b5d40_result_delayed_u0=1'h0;
reg		reg_00326d3c_result_delayed_u0=1'h0;
reg		reg_0f7fd2de_u0=1'h0;
reg		reg_27e96f4d_result_delayed_u0=1'h0;
reg		reg_57b67e1e_u0=1'h0;
reg		reg_2c075897_result_delayed_result_delayed_u0=1'h0;
reg		reg_6d65c4c8_u0=1'h0;
reg		reg_701b11b5_u0=1'h0;
reg		reg_7ff55f76_result_delayed_u0=1'h0;
reg		reg_6685c38c_result_delayed_u0=1'h0;
reg		reg_0edfde7a_result_delayed_result_delayed_u0=1'h0;
reg		reg_258519cc_result_delayed_u0=1'h0;
reg		reg_0c422d83_u0=1'h0;
reg		reg_6fbb03a9_result_delayed_u0=1'h0;
reg		reg_78fa2139_u0=1'h0;
reg		reg_0e4a778e_u0=1'h0;
reg		reg_00bce4e8_result_delayed_u0=1'h0;
reg		reg_56eb272e_u0=1'h0;
reg		reg_710c3541_result_delayed_u0=1'h0;
reg		reg_13e83e22_u0=1'h0;
reg		reg_2309bac6_u0=1'h0;
reg		reg_2eae6f7e_u0=1'h0;
reg		reg_2e62ff2a_result_delayed_u0=1'h0;
reg		reg_63ada2d0_result_delayed_u0=1'h0;
reg		reg_17d8460a_u0=1'h0;
reg		reg_63314f9f_result_delayed_u0=1'h0;
reg		reg_792a283d_result_delayed_u0=1'h0;
reg		reg_4ec17b1d_u0=1'h0;
reg		reg_74e3dda4_result_delayed_u0=1'h0;
reg		reg_6cf5c92b_u0=1'h0;
reg		reg_2cb89c91_result_delayed_u0=1'h0;
reg		reg_1a836fd8_result_delayed_u0=1'h0;
reg		reg_3e384fda_u0=1'h0;
reg		reg_5fd2d636_u0=1'h0;
reg		reg_09c6d144_result_delayed_u0=1'h0;
reg		reg_279d2f74_result_delayed_u0=1'h0;
reg		reg_3b4652ae_u0=1'h0;
reg		reg_52747b9c_u0=1'h0;
reg		reg_689d5d75_u0=1'h0;
reg		reg_00bce4e8_result_delayed_result_delayed_u0=1'h0;
reg		reg_6f7d9e94_u0=1'h0;
reg		reg_138117ea_result_delayed_u0=1'h0;
reg		reg_5acdfb21_u0=1'h0;
reg		reg_1de599bc_result_delayed_result_delayed_u0=1'h0;
reg		reg_030c675e_result_delayed_u0=1'h0;
reg		reg_437f3245_result_delayed_u0=1'h0;
reg		reg_63daa7a1_result_delayed_u0=1'h0;
reg		reg_258519cc_result_delayed_result_delayed_u0=1'h0;
reg		reg_158b107d_u0=1'h0;
reg		reg_5c74f06b_result_delayed_u0=1'h0;
reg		reg_54cc0137_u0=1'h0;
reg		reg_57713ae7_result_delayed_u0=1'h0;
reg		reg_0a0626a2_result_delayed_u0=1'h0;
reg		reg_36b55f4a_u0=1'h0;
reg		reg_05644f67_u0=1'h0;
reg		reg_25493747_u0=1'h0;
reg		reg_6741a229_result_delayed_u0=1'h0;
reg		reg_14e9d2f9_u0=1'h0;
reg		reg_7c5e48af_result_delayed_u0=1'h0;
reg		reg_47eb2b6a_result_delayed_u0=1'h0;
reg		reg_1de599bc_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_7c5e48af_result_delayed_result_delayed_u0=1'h0;
reg		reg_0bd3d5c5_u0=1'h0;
reg		reg_0e47a050_u0=1'h0;
reg		reg_76b494ad_u0=1'h0;
reg		reg_47f4e6ec_result_delayed_u0=1'h0;
reg		reg_792ef732_u0=1'h0;
reg		reg_678f3d92_u0=1'h0;
reg		reg_23499f80_result_delayed_u0=1'h0;
reg		reg_2309bac6_result_delayed_u0=1'h0;
reg		reg_2ca30e82_u0=1'h0;
reg		reg_58bcae9f_u0=1'h0;
reg		reg_701b11b5_result_delayed_u0=1'h0;
reg		reg_175ea576_u0=1'h0;
reg		reg_0cb5aa9c_u0=1'h0;
reg		reg_77dbf5f0_u0=1'h0;
reg		reg_5acdfb21_result_delayed_u0=1'h0;
reg		reg_3575e35b_u0=1'h0;
reg		reg_7c5e48af_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_18cb5efb_u0=1'h0;
reg		reg_59c65bf7_u0=1'h0;
reg		reg_701b11b5_result_delayed_result_delayed_u0=1'h0;
reg		reg_2f53bd66_u0=1'h0;
reg		reg_4cf96ace_u0=1'h0;
reg		reg_33167b6e_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_515acf62_u0=1'h0;
reg		reg_37bbd983_u0=1'h0;
reg		reg_640558fa_result_delayed_u0=1'h0;
reg		reg_7d614f5b_u0=1'h0;
reg		reg_78fa2139_result_delayed_u0=1'h0;
reg		reg_17699155_u0=1'h0;
reg		reg_5fd2d636_result_delayed_u0=1'h0;
reg		reg_09c6d144_result_delayed_result_delayed_u0=1'h0;
reg		reg_792a283d_result_delayed_result_delayed_u0=1'h0;
reg		reg_7dd4b39e_u0=1'h0;
reg		reg_2dac7bf9_u0=1'h0;
reg		reg_107844c4_result_delayed_result_delayed_u0=1'h0;
reg		reg_33b11310_result_delayed_u0=1'h0;
reg		reg_5aa7d6c8_result_delayed_u0=1'h0;
reg		reg_77047715_result_delayed_u0=1'h0;
reg		reg_03e66f15_result_delayed_u0=1'h0;
reg		reg_530b2d69_u0=1'h0;
reg		reg_0a611af4_result_delayed_u0=1'h0;
reg		reg_3e784e1c_result_delayed_result_delayed_u0=1'h0;
reg		reg_5fc6e1a0_u0=1'h0;
reg		reg_3b393219_result_delayed_u0=1'h0;
reg		reg_70cebea7_u0=1'h0;
reg		reg_31796710_u0=1'h0;
reg		reg_370ead64_u0=1'h0;
reg		reg_62f7fc9b_u0=1'h0;
reg		reg_05fe2b93_u0=1'h0;
reg		reg_01db913f_result_delayed_u0=1'h0;
reg		reg_3c118266_u0=1'h0;
reg		reg_32fe623a_result_delayed_u0=1'h0;
reg		reg_387e0416_result_delayed_u0=1'h0;
reg		reg_1dd4f50d_result_delayed_u0=1'h0;
reg		reg_64870a03_u0=1'h0;
reg		reg_7a88ee59_result_delayed_result_delayed_u0=1'h0;
reg		reg_485faada_u0=1'h0;
reg		reg_7c7216f8_u0=1'h0;
reg		reg_689528f4_result_delayed_result_delayed_u0=1'h0;
reg		and_delayed_u207=1'h0;
reg		reg_42afe023_u0=1'h0;
reg		reg_6fbb03a9_result_delayed_result_delayed_u0=1'h0;
reg		reg_0a611af4_result_delayed_result_delayed_u0=1'h0;
reg		reg_33b11310_result_delayed_result_delayed_u0=1'h0;
reg		reg_3d06bf89_u0=1'h0;
reg		reg_17fed16d_u0=1'h0;
reg		reg_3f347781_result_delayed_u0=1'h0;
wire		mux_u315;
wire		or_u895_u0;
reg		reg_279d2f74_result_delayed_result_delayed_u0=1'h0;
reg		reg_54cc0137_result_delayed_u0=1'h0;
reg		reg_27e96f4d_result_delayed_result_delayed_u0=1'h0;
reg		reg_57b67e1e_result_delayed_u0=1'h0;
reg		reg_355135b7_result_delayed_result_delayed_u0=1'h0;
reg		reg_1536340b_result_delayed_u0=1'h0;
reg		reg_3c99258f_result_delayed_u0=1'h0;
reg		reg_05fe2b93_result_delayed_u0=1'h0;
reg		reg_4b516dfb_u0=1'h0;
reg		reg_6e43fb69_result_delayed_u0=1'h0;
reg		reg_7c7f1881_result_delayed_u0=1'h0;
reg		reg_04854db4_result_delayed_u0=1'h0;
reg		reg_3e384fda_result_delayed_u0=1'h0;
reg		reg_09c6d144_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_3715a5a1_u0=1'h0;
reg		reg_33b11310_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_62f7fc9b_result_delayed_u0=1'h0;
reg		reg_54fa2642_u0=1'h0;
reg		reg_44204699_u0=1'h0;
reg		reg_03ce3977_u0=1'h0;
reg		reg_28399a83_u0=1'h0;
reg		reg_57713ae7_result_delayed_result_delayed_u0=1'h0;
reg		reg_2ecaeed5_result_delayed_result_delayed_u0=1'h0;
reg		reg_2a1c2b8c_result_delayed_u0=1'h0;
reg		reg_78fa2139_result_delayed_result_delayed_u0=1'h0;
reg		reg_7a88ee59_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_40adac30_result_delayed_result_delayed_u0=1'h0;
reg		reg_2dac7bf9_result_delayed_u0=1'h0;
reg		reg_5085924e_u0=1'h0;
reg		reg_6d657fae_u0=1'h0;
reg		reg_05074d01_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_18cb5efb_result_delayed_u0=1'h0;
reg		reg_77b9b56b_u0=1'h0;
reg		reg_7bc1bfcd_result_delayed_u0=1'h0;
reg		reg_0edfde7a_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_2c3cec3a_result_delayed_u0=1'h0;
reg		reg_5fc6e1a0_result_delayed_u0=1'h0;
reg		reg_107844c4_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_2349ca1b_result_delayed_u0=1'h0;
reg		reg_4d6a0c19_result_delayed_u0=1'h0;
reg		reg_546fd8be_result_delayed_u0=1'h0;
reg		reg_2c075897_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_57b67e1e_result_delayed_result_delayed_u0=1'h0;
reg		reg_429ea278_result_delayed_u0=1'h0;
reg		reg_711087ce_u0=1'h0;
reg		reg_2d3a4979_result_delayed_u0=1'h0;
reg		reg_5f584dbb_u0=1'h0;
reg		reg_35da391c_result_delayed_u0=1'h0;
reg		reg_258519cc_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_13e83e22_result_delayed_u0=1'h0;
reg		reg_43b7c159_u0=1'h0;
reg		reg_00326d3c_result_delayed_result_delayed_u0=1'h0;
reg		reg_1de599bc_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_71bdf9cc_result_delayed_u0=1'h0;
reg		reg_1a836fd8_result_delayed_result_delayed_u0=1'h0;
reg		reg_2ca30e82_result_delayed_u0=1'h0;
reg		reg_5b15db0b_result_delayed_u0=1'h0;
reg		reg_0a6e669d_result_delayed_u0=1'h0;
reg		reg_54cc0137_result_delayed_result_delayed_u0=1'h0;
reg		reg_2eae6f7e_result_delayed_u0=1'h0;
reg		reg_0fb3eac1_result_delayed_u0=1'h0;
reg		reg_5011c507_result_delayed_u0=1'h0;
reg		reg_32e22ff9_result_delayed_u0=1'h0;
reg		reg_43d5e336_result_delayed_u0=1'h0;
reg		reg_05286558_result_delayed_u0=1'h0;
reg		reg_14e9d2f9_result_delayed_u0=1'h0;
reg		reg_5d8c3e8b_u0=1'h0;
reg		reg_0bfe7f33_result_delayed_u0=1'h0;
reg		reg_05fe2b93_result_delayed_result_delayed_u0=1'h0;
reg		reg_03e66f15_result_delayed_result_delayed_u0=1'h0;
reg		reg_50917495_result_delayed_u0=1'h0;
reg		reg_770cdc1d_u0=1'h0;
reg		reg_258519cc_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_7b23ef69_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_09c6d144_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_5c72dd07_result_delayed_u0=1'h0;
reg		reg_77dbf5f0_result_delayed_u0=1'h0;
reg		reg_1536340b_result_delayed_result_delayed_u0=1'h0;
reg		reg_0304da20_result_delayed_result_delayed_u0=1'h0;
reg		reg_401b0405_result_delayed_u0=1'h0;
reg		reg_50917495_result_delayed_result_delayed_u0=1'h0;
reg		reg_682b29b0_result_delayed_u0=1'h0;
reg		reg_7a3ed379_result_delayed_u0=1'h0;
reg		reg_66095291_result_delayed_u0=1'h0;
reg		reg_7ec4fde8_u0=1'h0;
reg		reg_0e12093d_u0=1'h0;
reg		reg_689528f4_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_0c422d83_result_delayed_u0=1'h0;
reg		reg_31796710_result_delayed_u0=1'h0;
reg		reg_062c6117_u0=1'h0;
reg		reg_41025437_result_delayed_u0=1'h0;
wire		and_u3151_u0;
reg		reg_5fd2d636_result_delayed_result_delayed_u0=1'h0;
reg		reg_23b56b6a_result_delayed_u0=1'h0;
reg		reg_318c1131_result_delayed_u0=1'h0;
reg		reg_638aaf04_result_delayed_u0=1'h0;
reg		reg_74c8f38e_u0=1'h0;
reg		reg_638aaf04_result_delayed_result_delayed_u0=1'h0;
reg		reg_41bcb2f2_u0=1'h0;
reg		reg_2a1f0d51_u0=1'h0;
reg		reg_1ca67dbd_result_delayed_u0=1'h0;
reg		reg_63daa7a1_result_delayed_result_delayed_u0=1'h0;
reg		reg_05fa154c_result_delayed_result_delayed_u0=1'h0;
reg		reg_37bbd983_result_delayed_u0=1'h0;
reg		reg_6741a229_result_delayed_result_delayed_u0=1'h0;
reg		reg_6741a229_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_1db07eea_u0=1'h0;
reg		reg_0afd59a6_u0=1'h0;
reg		reg_0e12093d_result_delayed_u0=1'h0;
reg		reg_15387666_u0=1'h0;
reg		reg_5780a32a_result_delayed_u0=1'h0;
reg		reg_3ac681a6_u0=1'h0;
reg		reg_792a283d_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_64870a03_result_delayed_u0=1'h0;
reg		reg_678f3d92_result_delayed_u0=1'h0;
reg		reg_387e0416_result_delayed_result_delayed_u0=1'h0;
reg		reg_049d2474_result_delayed_u0=1'h0;
reg		reg_711087ce_result_delayed_u0=1'h0;
reg		reg_3b4c4b37_result_delayed_u0=1'h0;
reg		reg_33b11310_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_20570b20_u0=1'h0;
reg		reg_37bbd983_result_delayed_result_delayed_u0=1'h0;
reg		reg_2a1f0d51_result_delayed_u0=1'h0;
reg		reg_55180568_result_delayed_u0=1'h0;
reg		reg_70cebea7_result_delayed_u0=1'h0;
reg		reg_297a657a_result_delayed_u0=1'h0;
reg		reg_5aa7d6c8_result_delayed_result_delayed_u0=1'h0;
reg		reg_47f4e6ec_result_delayed_result_delayed_u0=1'h0;
reg		reg_1b8047bd_result_delayed_u0=1'h0;
reg		reg_7f7d622f_result_delayed_u0=1'h0;
reg		reg_5011c507_result_delayed_result_delayed_u0=1'h0;
reg		reg_539db809_u0=1'h0;
reg		reg_0bfe7f33_result_delayed_result_delayed_u0=1'h0;
reg		reg_40e76b7d_u0=1'h0;
reg		reg_40d160ea_result_delayed_u0=1'h0;
reg		reg_7217fecc_result_delayed_u0=1'h0;
reg		reg_4e012e31_result_delayed_u0=1'h0;
reg		reg_7ff55f76_result_delayed_result_delayed_u0=1'h0;
reg		reg_6d5cb91c_result_delayed_u0=1'h0;
reg		reg_5f68d729_result_delayed_u0=1'h0;
reg		reg_3715a5a1_result_delayed_u0=1'h0;
reg		reg_41025437_result_delayed_result_delayed_u0=1'h0;
reg		reg_6109ede1_result_delayed_u0=1'h0;
reg		reg_4a292b3c_result_delayed_u0=1'h0;
reg		reg_7ec4fde8_result_delayed_u0=1'h0;
reg		reg_378e778c_result_delayed_u0=1'h0;
reg		reg_64fa00de_result_delayed_result_delayed_u0=1'h0;
reg		reg_0e47a050_result_delayed_u0=1'h0;
reg		reg_17e75387_result_delayed_u0=1'h0;
reg		reg_3d4ff93c_result_delayed_u0=1'h0;
reg		reg_15387666_result_delayed_u0=1'h0;
reg		reg_12289738_result_delayed_u0=1'h0;
reg		reg_74e3dda4_result_delayed_result_delayed_u0=1'h0;
reg		reg_4b39e741_result_delayed_u0=1'h0;
reg		reg_54826c24_result_delayed_u0=1'h0;
reg		reg_297a657a_result_delayed_result_delayed_u0=1'h0;
reg		reg_6806d06c_result_delayed_u0=1'h0;
reg		reg_0c3478e6_result_delayed_result_delayed_u0=1'h0;
reg		reg_1536c80b_result_delayed_u0=1'h0;
reg		reg_7a51229e_result_delayed_u0=1'h0;
reg		reg_6dc4bd1b_result_delayed_u0=1'h0;
reg		reg_43039f69_result_delayed_result_delayed_u0=1'h0;
reg		reg_5780a32a_result_delayed_result_delayed_u0=1'h0;
reg		reg_29782e98_u0=1'h0;
reg		reg_536a7781_result_delayed_u0=1'h0;
reg		reg_32a6867b_result_delayed_result_delayed_u0=1'h0;
reg		reg_683a6054_result_delayed_u0=1'h0;
reg		reg_58bcae9f_result_delayed_u0=1'h0;
reg		reg_7d614f5b_result_delayed_u0=1'h0;
reg		reg_57b67e1e_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_4cf96ace_result_delayed_u0=1'h0;
reg		reg_35ff7cc6_result_delayed_u0=1'h0;
reg		and_delayed_u208_u0=1'h0;
wire		or_u896_u0;
reg		reg_77b9b56b_result_delayed_u0=1'h0;
wire		or_u897_u0;
wire		and_u3152_u0;
wire		and_u3153_u0;
wire		or_u898_u0;
wire		mux_u316_u0;
reg		reg_58165587_u0=1'h0;
wire		or_u899_u0;
wire	[31:0]	mux_u317_u0;
wire		or_u900_u0;
reg		reg_31cf41da_u0=1'h0;
wire		or_u901_u0;
wire		or_u902_u0;
reg		and_delayed_u209_u0=1'h0;
wire		and_u3154_u0;
wire		and_u3155_u0;
wire		or_u903_u0;
reg		and_delayed_u210_u0=1'h0;
wire signed	[31:0]	equals_u166_a_signed;
wire signed	[31:0]	equals_u166_b_signed;
wire		equals_u166;
wire		and_u3156_u0;
wire		not_u530_u0;
wire		and_u3157_u0;
wire		and_u3158_u0;
wire		not_u531_u0;
wire		and_u3159_u0;
wire		lessThan_u75;
wire signed	[31:0]	lessThan_u75_a_signed;
wire signed	[31:0]	lessThan_u75_b_signed;
wire		and_u3160_u0;
wire		and_u3161_u0;
wire		not_u532_u0;
wire		and_u3162_u0;
wire		and_u3163_u0;
wire		not_u533_u0;
wire	[31:0]	add;
wire		and_u3164_u0;
wire	[15:0]	simplePinWrite_u468;
wire	[15:0]	simplePinWrite_u469;
wire		simplePinWrite_u470;
wire	[31:0]	add_u374;
reg	[15:0]	syncEnable_u550=16'h0;
wire		and_u3165_u0;
reg		reg_0de2a3c0_u0=1'h0;
reg		and_delayed_u211_u0=1'h0;
wire	[15:0]	mux_u318_u0;
reg	[15:0]	syncEnable_u551_u0=16'h0;
wire		and_u3166_u0;
reg		reg_0498419c_u0=1'h0;
wire	[15:0]	mux_u319_u0;
wire	[31:0]	mux_u320_u0;
reg	[31:0]	syncEnable_u552_u0=32'h0;
reg	[15:0]	syncEnable_u553_u0=16'h0;
wire		and_u3167_u0;
reg		and_delayed_u212_u0=1'h0;
wire		and_u3168_u0;
reg		reg_490a59eb_u0=1'h0;
wire	[15:0]	mux_u321_u0;
wire	[31:0]	mux_u322_u0;
reg		reg_5602ca0c_u0=1'h0;
wire		and_u3169_u0;
reg	[15:0]	syncEnable_u554_u0=16'h0;
reg	[31:0]	syncEnable_u555_u0=32'h0;
wire		and_u3170_u0;
wire	[15:0]	mux_u323_u0;
wire		and_u3171_u0;
reg	[31:0]	syncEnable_u556_u0=32'h0;
wire	[31:0]	mux_u324_u0;
reg		reg_7e9a4e4d_u0=1'h0;
reg		and_delayed_u213_u0=1'h0;
wire		and_u3172_u0;
reg	[15:0]	syncEnable_u557_u0=16'h0;
reg	[15:0]	latch_3dab8262_reg=16'h0;
wire	[15:0]	latch_3dab8262_out;
wire		mux_u325_u0;
wire		or_u904_u0;
wire		or_u905_u0;
wire		mux_u326_u0;
reg	[31:0]	latch_182feb1c_reg=32'h0;
wire	[31:0]	latch_182feb1c_out;
wire	[31:0]	mux_u327_u0;
wire		or_u906_u0;
wire	[31:0]	mux_u328_u0;
wire		or_u907_u0;
reg		block_GO_delayed_u10=1'h0;
reg	[31:0]	fbReg_temp_fsmOldState_resized_LH1_xy_6_u0=32'h0;
wire	[15:0]	mux_u329_u0;
wire	[31:0]	mux_u330_u0;
reg	[15:0]	fbReg_Out1Portvalue_u3=16'h0;
reg		syncEnable_u558_u0=1'h0;
reg		loopControl_u7=1'h0;
wire		or_u908_u0;
wire	[31:0]	mux_u331_u0;
wire		or_u909_u0;
reg		reg_687233e3_u0=1'h0;
wire		or_u910_u0;
wire		mux_u332_u0;
wire		or_u911_u0;
wire		mux_u333_u0;
wire		or_u912_u0;
reg		reg_687233e3_result_delayed_u0=1'h0;
wire	[31:0]	mux_u334_u0;
wire		or_u913_u0;
assign and_u3140_u0=or_u908_u0&or_u908_u0;
assign lessThan_a_unsigned=port_008a440f_;
assign lessThan_b_unsigned=16'h100;
assign lessThan=lessThan_a_unsigned<lessThan_b_unsigned;
assign equals_a_unsigned=port_008a440f_;
assign equals_b_unsigned=16'h100;
assign equals=equals_a_unsigned==equals_b_unsigned;
assign lessThan_u74_a_unsigned=port_1ba874b3_;
assign lessThan_u74_b_unsigned=16'h2;
assign lessThan_u74=lessThan_u74_a_unsigned<lessThan_u74_b_unsigned;
assign andOp=equals&lessThan_u74;
assign equals_u164_a_unsigned=port_1ba874b3_;
assign equals_u164_b_unsigned=16'h2;
assign equals_u164=equals_u164_a_unsigned==equals_u164_b_unsigned;
assign equals_u165_a_signed={31'b0, port_0a81f2c6_};
assign equals_u165_b_signed=32'h0;
assign equals_u165=equals_u165_a_signed==equals_u165_b_signed;
assign not_u526_u0=~equals_u165;
assign and_u3141_u0=and_u3140_u0&not_u526_u0;
assign and_u3142_u0=and_u3140_u0&equals_u165;
assign andOp_u173=lessThan&port_58303e5a_;
assign and_u3143_u0=and_u3155_u0&not_u527_u0;
assign and_u3144_u0=and_u3155_u0&andOp_u173;
assign not_u527_u0=~andOp_u173;
assign simplePinWrite=and_u3153_u0&{1{and_u3153_u0}};
assign and_u3145_u0=and_u3152_u0&andOp;
assign not_u528_u0=~andOp;
assign and_u3146_u0=and_u3152_u0&not_u528_u0;
assign simplePinWrite_u466=and_u3150_u0&{1{and_u3150_u0}};
assign and_u3147_u0=and_u3151_u0&equals_u164;
assign not_u529_u0=~equals_u164;
assign and_u3148_u0=and_u3151_u0&not_u529_u0;
assign simplePinWrite_u467=and_u3149_u0&{1{and_u3149_u0}};
assign and_u3149_u0=and_u3147_u0&and_u3151_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_297a657a_u0<=1'h0;
else reg_297a657a_u0<=reg_258519cc_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_378e778c_u0<=1'h0;
else reg_378e778c_u0<=reg_79b769ec_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_50917495_u0<=1'h0;
else reg_50917495_u0<=reg_342c7170_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_05074d01_u0<=1'h0;
else reg_05074d01_u0<=reg_3ac681a6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2c3cec3a_u0<=1'h0;
else reg_2c3cec3a_u0<=reg_77047715_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7bc1bfcd_u0<=1'h0;
else reg_7bc1bfcd_u0<=reg_05c10dfa_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_77047715_u0<=1'h0;
else reg_77047715_u0<=reg_18cb5efb_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6fbb03a9_u0<=1'h0;
else reg_6fbb03a9_u0<=reg_2139e56a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_401b0405_u0<=1'h0;
else reg_401b0405_u0<=reg_5085924e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5b15db0b_u0<=1'h0;
else reg_5b15db0b_u0<=reg_281f24ad_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5c74f06b_u0<=1'h0;
else reg_5c74f06b_u0<=reg_1ab96b28_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2ecaeed5_u0<=1'h0;
else reg_2ecaeed5_u0<=reg_6e8b025a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_64fa00de_u0<=1'h0;
else reg_64fa00de_u0<=reg_324e3a7d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_65acfd8b_u0<=1'h0;
else reg_65acfd8b_u0<=reg_57b67e1e_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2cb89c91_u0<=1'h0;
else reg_2cb89c91_u0<=reg_1a7a9643_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4e012e31_u0<=1'h0;
else reg_4e012e31_u0<=reg_175ea576_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_324e3a7d_u0<=1'h0;
else reg_324e3a7d_u0<=reg_429ea278_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_324e3a7d_result_delayed_u0<=1'h0;
else reg_324e3a7d_result_delayed_u0<=reg_324e3a7d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1a7a9643_u0<=1'h0;
else reg_1a7a9643_u0<=reg_7e56828a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_40d160ea_u0<=1'h0;
else reg_40d160ea_u0<=reg_4e70c2f7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_05c10dfa_u0<=1'h0;
else reg_05c10dfa_u0<=reg_5e96aee9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_357b5d40_u0<=1'h0;
else reg_357b5d40_u0<=reg_60f891d5_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1b8047bd_u0<=1'h0;
else reg_1b8047bd_u0<=reg_00326d3c_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6d5cb91c_u0<=1'h0;
else reg_6d5cb91c_u0<=reg_6b6d7306_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5f68d729_u0<=1'h0;
else reg_5f68d729_u0<=reg_4d6a0c19_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2d3a4979_u0<=1'h0;
else reg_2d3a4979_u0<=reg_14fc4001_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_258519cc_u0<=1'h0;
else reg_258519cc_u0<=reg_0edfde7a_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7b23ef69_u0<=1'h0;
else reg_7b23ef69_u0<=reg_52d98a27_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4e9c06d0_u0<=1'h0;
else reg_4e9c06d0_u0<=reg_01aa19f9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_710c3541_u0<=1'h0;
else reg_710c3541_u0<=reg_3575e35b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6e5ada14_u0<=1'h0;
else reg_6e5ada14_u0<=reg_638aaf04_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_030c675e_u0<=1'h0;
else reg_030c675e_u0<=reg_678f3d92_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2139e56a_u0<=1'h0;
else reg_2139e56a_u0<=reg_04854db4_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01aa19f9_u0<=1'h0;
else reg_01aa19f9_u0<=reg_1b57bf2f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00bce4e8_u0<=1'h0;
else reg_00bce4e8_u0<=reg_65acfd8b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1de599bc_u0<=1'h0;
else reg_1de599bc_u0<=reg_7c7216f8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_79b769ec_u0<=1'h0;
else reg_79b769ec_u0<=reg_6e5ada14_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_17e75387_u0<=1'h0;
else reg_17e75387_u0<=reg_0cb5aa9c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_689528f4_u0<=1'h0;
else reg_689528f4_u0<=reg_1f49a7e5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3e784e1c_u0<=1'h0;
else reg_3e784e1c_u0<=reg_0c3478e6_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_387e0416_u0<=1'h0;
else reg_387e0416_u0<=reg_0f7fd2de_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_43039f69_u0<=1'h0;
else reg_43039f69_u0<=reg_74e3dda4_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6806d06c_u0<=1'h0;
else reg_6806d06c_u0<=reg_2309bac6_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6b6d7306_u0<=1'h0;
else reg_6b6d7306_u0<=reg_3f347781_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_138117ea_u0<=1'h0;
else reg_138117ea_u0<=reg_2f53bd66_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_683a6054_u0<=1'h0;
else reg_683a6054_u0<=reg_5f095be9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5aa7d6c8_u0<=1'h0;
else reg_5aa7d6c8_u0<=reg_0e47a050_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_05286558_u0<=1'h0;
else reg_05286558_u0<=reg_49dd354a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_55180568_u0<=1'h0;
else reg_55180568_u0<=reg_2bfa4eac_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_71bdf9cc_u0<=1'h0;
else reg_71bdf9cc_u0<=reg_485faada_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_79b769ec_result_delayed_u0<=1'h0;
else reg_79b769ec_result_delayed_u0<=reg_79b769ec_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3d4ff93c_u0<=1'h0;
else reg_3d4ff93c_u0<=reg_49f0052b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1b57bf2f_u0<=1'h0;
else reg_1b57bf2f_u0<=reg_43d5e336_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_33167b6e_u0<=1'h0;
else reg_33167b6e_u0<=reg_7a88ee59_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4b39e741_u0<=1'h0;
else reg_4b39e741_u0<=reg_4b516dfb_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_63daa7a1_u0<=1'h0;
else reg_63daa7a1_u0<=reg_3c8b940e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3b4c4b37_u0<=1'h0;
else reg_3b4c4b37_u0<=reg_40d160ea_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5e96aee9_u0<=1'h0;
else reg_5e96aee9_u0<=reg_0e4a778e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_47eb2b6a_u0<=1'h0;
else reg_47eb2b6a_u0<=reg_3212b28a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_09c6d144_u0<=1'h0;
else reg_09c6d144_u0<=reg_437f3245_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7ff55f76_u0<=1'h0;
else reg_7ff55f76_u0<=reg_43b7c159_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3c8b940e_u0<=1'h0;
else reg_3c8b940e_u0<=reg_6a06c71e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4e70c2f7_u0<=1'h0;
else reg_4e70c2f7_u0<=reg_370ead64_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6e5ada14_result_delayed_u0<=1'h0;
else reg_6e5ada14_result_delayed_u0<=reg_6e5ada14_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3e784e1c_result_delayed_u0<=1'h0;
else reg_3e784e1c_result_delayed_u0<=reg_3e784e1c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_638aaf04_u0<=1'h0;
else reg_638aaf04_u0<=reg_76b494ad_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2c075897_u0<=1'h0;
else reg_2c075897_u0<=reg_63c2bf6e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0a611af4_u0<=1'h0;
else reg_0a611af4_u0<=reg_3b4652ae_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_49dd354a_u0<=1'h0;
else reg_49dd354a_u0<=reg_401b0405_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3212b28a_u0<=1'h0;
else reg_3212b28a_u0<=reg_2c075897_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_66095291_u0<=1'h0;
else reg_66095291_u0<=reg_2f7313b9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_40adac30_u0<=1'h0;
else reg_40adac30_u0<=reg_5f7ee655_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_33b11310_u0<=1'h0;
else reg_33b11310_u0<=reg_6685c38c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_27e96f4d_u0<=1'h0;
else reg_27e96f4d_u0<=reg_792ef732_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0a0626a2_u0<=1'h0;
else reg_0a0626a2_u0<=reg_50917495_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0edfde7a_u0<=1'h0;
else reg_0edfde7a_u0<=reg_5cd43dad_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_54826c24_u0<=1'h0;
else reg_54826c24_u0<=reg_10dd85da_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_43039f69_result_delayed_u0<=1'h0;
else reg_43039f69_result_delayed_u0<=reg_43039f69_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5780a32a_u0<=1'h0;
else reg_5780a32a_u0<=reg_1de599bc_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_63c2bf6e_u0<=1'h0;
else reg_63c2bf6e_u0<=reg_2dac7bf9_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1f49a7e5_u0<=1'h0;
else reg_1f49a7e5_u0<=reg_6d65c4c8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_63314f9f_u0<=1'h0;
else reg_63314f9f_u0<=reg_0afd59a6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_281f24ad_u0<=1'h0;
else reg_281f24ad_u0<=reg_2349ca1b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3212b28a_result_delayed_u0<=1'h0;
else reg_3212b28a_result_delayed_u0<=reg_3212b28a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3f347781_u0<=1'h0;
else reg_3f347781_u0<=reg_29259ddf_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_05fa154c_u0<=1'h0;
else reg_05fa154c_u0<=reg_4cf96ace_result_delayed_u0;
end
assign and_u3150_u0=and_u3145_u0&and_u3152_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2139e56a_result_delayed_u0<=1'h0;
else reg_2139e56a_result_delayed_u0<=reg_2139e56a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_107844c4_u0<=1'h0;
else reg_107844c4_u0<=reg_3e384fda_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_318c1131_u0<=1'h0;
else reg_318c1131_u0<=reg_31796710_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_689528f4_result_delayed_u0<=1'h0;
else reg_689528f4_result_delayed_u0<=reg_689528f4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_32fe623a_u0<=1'h0;
else reg_32fe623a_u0<=reg_2d3a4979_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_69fad53c_u0<=1'h0;
else reg_69fad53c_u0<=reg_6cf5c92b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_35da391c_u0<=1'h0;
else reg_35da391c_u0<=reg_5fc6e1a0_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_23499f80_u0<=1'h0;
else reg_23499f80_u0<=reg_75b844ca_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2f7313b9_u0<=1'h0;
else reg_2f7313b9_u0<=reg_689528f4_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2ecaeed5_result_delayed_u0<=1'h0;
else reg_2ecaeed5_result_delayed_u0<=reg_2ecaeed5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_107844c4_result_delayed_u0<=1'h0;
else reg_107844c4_result_delayed_u0<=reg_107844c4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0bfe7f33_u0<=1'h0;
else reg_0bfe7f33_u0<=reg_69fad53c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a51229e_u0<=1'h0;
else reg_7a51229e_u0<=reg_7c7f1881_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_33167b6e_result_delayed_u0<=1'h0;
else reg_33167b6e_result_delayed_u0<=reg_33167b6e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6e8b025a_u0<=1'h0;
else reg_6e8b025a_u0<=reg_5c74f06b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_546fd8be_u0<=1'h0;
else reg_546fd8be_u0<=reg_6fbb03a9_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a88ee59_u0<=1'h0;
else reg_7a88ee59_u0<=reg_6fc41285_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0c3478e6_u0<=1'h0;
else reg_0c3478e6_u0<=reg_64870a03_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1de599bc_result_delayed_u0<=1'h0;
else reg_1de599bc_result_delayed_u0<=reg_1de599bc_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_05074d01_result_delayed_u0<=1'h0;
else reg_05074d01_result_delayed_u0<=reg_05074d01_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1dd4f50d_u0<=1'h0;
else reg_1dd4f50d_u0<=reg_5eccd3e3_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_49f0052b_u0<=1'h0;
else reg_49f0052b_u0<=reg_3622ef46_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7217fecc_u0<=1'h0;
else reg_7217fecc_u0<=reg_5fd2d636_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7e56828a_u0<=1'h0;
else reg_7e56828a_u0<=reg_6d657fae_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_32a6867b_u0<=1'h0;
else reg_32a6867b_u0<=reg_1db07eea_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6dc4bd1b_u0<=1'h0;
else reg_6dc4bd1b_u0<=reg_03ce3977_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_23b56b6a_u0<=1'h0;
else reg_23b56b6a_u0<=reg_4b39e741_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0edfde7a_result_delayed_u0<=1'h0;
else reg_0edfde7a_result_delayed_u0<=reg_0edfde7a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5f095be9_u0<=1'h0;
else reg_5f095be9_u0<=reg_357b5d40_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_43d5e336_u0<=1'h0;
else reg_43d5e336_u0<=reg_0fb3eac1_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_64fa00de_result_delayed_u0<=1'h0;
else reg_64fa00de_result_delayed_u0<=reg_64fa00de_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01db913f_u0<=1'h0;
else reg_01db913f_u0<=reg_63ada2d0_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_355135b7_u0<=1'h0;
else reg_355135b7_u0<=reg_640558fa_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_429ea278_u0<=1'h0;
else reg_429ea278_u0<=reg_05fe2b93_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6109ede1_u0<=1'h0;
else reg_6109ede1_u0<=reg_1e58db1f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_049d2474_u0<=1'h0;
else reg_049d2474_u0<=reg_0319ee54_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_279d2f74_u0<=1'h0;
else reg_279d2f74_u0<=reg_6c0ed978_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_536a7781_u0<=1'h0;
else reg_536a7781_u0<=reg_25493747_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7c5e48af_u0<=1'h0;
else reg_7c5e48af_u0<=reg_41bcb2f2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_355135b7_result_delayed_u0<=1'h0;
else reg_355135b7_result_delayed_u0<=reg_355135b7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_03e66f15_u0<=1'h0;
else reg_03e66f15_u0<=reg_5a95fe6b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0a6e669d_u0<=1'h0;
else reg_0a6e669d_u0<=reg_279d2f74_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_29259ddf_u0<=1'h0;
else reg_29259ddf_u0<=reg_56eb272e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_14fc4001_u0<=1'h0;
else reg_14fc4001_u0<=reg_1dd4f50d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7c7f1881_u0<=1'h0;
else reg_7c7f1881_u0<=reg_05074d01_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5a95fe6b_u0<=1'h0;
else reg_5a95fe6b_u0<=reg_158b107d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_52d98a27_u0<=1'h0;
else reg_52d98a27_u0<=reg_530b2d69_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_640558fa_u0<=1'h0;
else reg_640558fa_u0<=reg_00bce4e8_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_05c10dfa_result_delayed_u0<=1'h0;
else reg_05c10dfa_result_delayed_u0<=reg_05c10dfa_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7b23ef69_result_delayed_u0<=1'h0;
else reg_7b23ef69_result_delayed_u0<=reg_7b23ef69_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_10dd85da_u0<=1'h0;
else reg_10dd85da_u0<=reg_5aa7d6c8_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6685c38c_u0<=1'h0;
else reg_6685c38c_u0<=and_delayed_u207;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00326d3c_u0<=1'h0;
else reg_00326d3c_u0<=reg_378e778c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_65acfd8b_result_delayed_u0<=1'h0;
else reg_65acfd8b_result_delayed_u0<=reg_65acfd8b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_12289738_u0<=1'h0;
else reg_12289738_u0<=reg_74c8f38e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_05fa154c_result_delayed_u0<=1'h0;
else reg_05fa154c_result_delayed_u0<=reg_05fa154c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4a292b3c_u0<=1'h0;
else reg_4a292b3c_u0<=reg_47eb2b6a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5011c507_u0<=1'h0;
else reg_5011c507_u0<=reg_52747b9c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3c99258f_u0<=1'h0;
else reg_3c99258f_u0<=reg_7c5e48af_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_792a283d_u0<=1'h0;
else reg_792a283d_u0<=reg_4e9c06d0_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6a06c71e_u0<=1'h0;
else reg_6a06c71e_u0<=reg_7dd4b39e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0c3478e6_result_delayed_u0<=1'h0;
else reg_0c3478e6_result_delayed_u0<=reg_0c3478e6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_47f4e6ec_u0<=1'h0;
else reg_47f4e6ec_u0<=reg_6741a229_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_32e22ff9_u0<=1'h0;
else reg_32e22ff9_u0<=reg_47b1c63c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1ca67dbd_u0<=1'h0;
else reg_1ca67dbd_u0<=reg_5b15db0b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3b393219_u0<=1'h0;
else reg_3b393219_u0<=reg_70cebea7_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0304da20_u0<=1'h0;
else reg_0304da20_u0<=reg_57713ae7_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_40adac30_result_delayed_u0<=1'h0;
else reg_40adac30_result_delayed_u0<=reg_40adac30_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6e43fb69_u0<=1'h0;
else reg_6e43fb69_u0<=reg_261ccf7a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5f7ee655_u0<=1'h0;
else reg_5f7ee655_u0<=reg_3bc4d242_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0304da20_result_delayed_u0<=1'h0;
else reg_0304da20_result_delayed_u0<=reg_0304da20_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_60f891d5_u0<=1'h0;
else reg_60f891d5_u0<=reg_17fed16d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5eccd3e3_u0<=1'h0;
else reg_5eccd3e3_u0<=reg_701b11b5_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_04854db4_u0<=1'h0;
else reg_04854db4_u0<=reg_17699155_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6b6d7306_result_delayed_u0<=1'h0;
else reg_6b6d7306_result_delayed_u0<=reg_6b6d7306_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_41025437_u0<=1'h0;
else reg_41025437_u0<=reg_66095291_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_35ff7cc6_u0<=1'h0;
else reg_35ff7cc6_u0<=reg_32fe623a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_437f3245_u0<=1'h0;
else reg_437f3245_u0<=reg_0e12093d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1536c80b_u0<=1'h0;
else reg_1536c80b_u0<=reg_7e0ad75d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1536340b_u0<=1'h0;
else reg_1536340b_u0<=reg_17d8460a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_33167b6e_result_delayed_result_delayed_u0<=1'h0;
else reg_33167b6e_result_delayed_result_delayed_u0<=reg_33167b6e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6fc41285_u0<=1'h0;
else reg_6fc41285_u0<=reg_11d4a896_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_11d4a896_u0<=1'h0;
else reg_11d4a896_u0<=reg_2dbd2c2b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_32a6867b_result_delayed_u0<=1'h0;
else reg_32a6867b_result_delayed_u0<=reg_32a6867b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4e9c06d0_result_delayed_u0<=1'h0;
else reg_4e9c06d0_result_delayed_u0<=reg_4e9c06d0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1e58db1f_u0<=1'h0;
else reg_1e58db1f_u0<=reg_27e96f4d_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_74e3dda4_u0<=1'h0;
else reg_74e3dda4_u0<=reg_0a0626a2_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a3ed379_u0<=1'h0;
else reg_7a3ed379_u0<=reg_33167b6e_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2e62ff2a_u0<=1'h0;
else reg_2e62ff2a_u0<=reg_4f8202d0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a88ee59_result_delayed_u0<=1'h0;
else reg_7a88ee59_result_delayed_u0<=reg_7a88ee59_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_05074d01_result_delayed_result_delayed_u0<=1'h0;
else reg_05074d01_result_delayed_result_delayed_u0<=reg_05074d01_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0319ee54_u0<=1'h0;
else reg_0319ee54_u0<=reg_2e62ff2a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4f8202d0_u0<=1'h0;
else reg_4f8202d0_u0<=reg_15387666_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2349ca1b_u0<=1'h0;
else reg_2349ca1b_u0<=reg_7d614f5b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7f7d622f_u0<=1'h0;
else reg_7f7d622f_u0<=reg_2cb89c91_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6e8b025a_result_delayed_u0<=1'h0;
else reg_6e8b025a_result_delayed_u0<=reg_6e8b025a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2bfa4eac_u0<=1'h0;
else reg_2bfa4eac_u0<=reg_6812ad6d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7e0ad75d_u0<=1'h0;
else reg_7e0ad75d_u0<=reg_09c6d144_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7b23ef69_result_delayed_result_delayed_u0<=1'h0;
else reg_7b23ef69_result_delayed_result_delayed_u0<=reg_7b23ef69_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1a836fd8_u0<=1'h0;
else reg_1a836fd8_u0<=reg_28399a83_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_342c7170_u0<=1'h0;
else reg_342c7170_u0<=reg_62f7fc9b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_69fad53c_result_delayed_u0<=1'h0;
else reg_69fad53c_result_delayed_u0<=reg_69fad53c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3622ef46_u0<=1'h0;
else reg_3622ef46_u0<=reg_5d8c3e8b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_261ccf7a_u0<=1'h0;
else reg_261ccf7a_u0<=reg_0bd3d5c5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6741a229_u0<=1'h0;
else reg_6741a229_u0<=reg_36b55f4a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_29259ddf_result_delayed_u0<=1'h0;
else reg_29259ddf_result_delayed_u0<=reg_29259ddf_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0fb3eac1_u0<=1'h0;
else reg_0fb3eac1_u0<=reg_387e0416_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_75b844ca_u0<=1'h0;
else reg_75b844ca_u0<=reg_35da391c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4d6a0c19_u0<=1'h0;
else reg_4d6a0c19_u0<=reg_710c3541_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_281f24ad_result_delayed_u0<=1'h0;
else reg_281f24ad_result_delayed_u0<=reg_281f24ad_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5c72dd07_u0<=1'h0;
else reg_5c72dd07_u0<=reg_7106847e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2c075897_result_delayed_u0<=1'h0;
else reg_2c075897_result_delayed_u0<=reg_2c075897_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6c0ed978_u0<=1'h0;
else reg_6c0ed978_u0<=reg_689d5d75_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7106847e_u0<=1'h0;
else reg_7106847e_u0<=reg_2a1c2b8c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5cd43dad_u0<=1'h0;
else reg_5cd43dad_u0<=reg_1b8047bd_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_63ada2d0_u0<=1'h0;
else reg_63ada2d0_u0<=reg_59c65bf7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6812ad6d_u0<=1'h0;
else reg_6812ad6d_u0<=reg_05644f67_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_14fc4001_result_delayed_u0<=1'h0;
else reg_14fc4001_result_delayed_u0<=reg_14fc4001_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3bc4d242_u0<=1'h0;
else reg_3bc4d242_u0<=reg_5c72dd07_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_47b1c63c_u0<=1'h0;
else reg_47b1c63c_u0<=reg_23b56b6a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2a1c2b8c_u0<=1'h0;
else reg_2a1c2b8c_u0<=reg_539db809_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1ab96b28_u0<=1'h0;
else reg_1ab96b28_u0<=reg_2eae6f7e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_60f891d5_result_delayed_u0<=1'h0;
else reg_60f891d5_result_delayed_u0<=reg_60f891d5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_57713ae7_u0<=1'h0;
else reg_57713ae7_u0<=reg_5acdfb21_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2dbd2c2b_u0<=1'h0;
else reg_2dbd2c2b_u0<=reg_2ca30e82_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_682b29b0_u0<=1'h0;
else reg_682b29b0_u0<=reg_63314f9f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_357b5d40_result_delayed_u0<=1'h0;
else reg_357b5d40_result_delayed_u0<=reg_357b5d40_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00326d3c_result_delayed_u0<=1'h0;
else reg_00326d3c_result_delayed_u0<=reg_00326d3c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0f7fd2de_u0<=1'h0;
else reg_0f7fd2de_u0<=reg_47f4e6ec_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_27e96f4d_result_delayed_u0<=1'h0;
else reg_27e96f4d_result_delayed_u0<=reg_27e96f4d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_57b67e1e_u0<=1'h0;
else reg_57b67e1e_u0<=reg_2ecaeed5_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2c075897_result_delayed_result_delayed_u0<=1'h0;
else reg_2c075897_result_delayed_result_delayed_u0<=reg_2c075897_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6d65c4c8_u0<=1'h0;
else reg_6d65c4c8_u0<=reg_54fa2642_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_701b11b5_u0<=1'h0;
else reg_701b11b5_u0<=reg_58bcae9f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7ff55f76_result_delayed_u0<=1'h0;
else reg_7ff55f76_result_delayed_u0<=reg_7ff55f76_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6685c38c_result_delayed_u0<=1'h0;
else reg_6685c38c_result_delayed_u0<=reg_6685c38c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0edfde7a_result_delayed_result_delayed_u0<=1'h0;
else reg_0edfde7a_result_delayed_result_delayed_u0<=reg_0edfde7a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_258519cc_result_delayed_u0<=1'h0;
else reg_258519cc_result_delayed_u0<=reg_258519cc_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0c422d83_u0<=1'h0;
else reg_0c422d83_u0<=reg_14e9d2f9_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6fbb03a9_result_delayed_u0<=1'h0;
else reg_6fbb03a9_result_delayed_u0<=reg_6fbb03a9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_78fa2139_u0<=1'h0;
else reg_78fa2139_u0<=reg_42afe023_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0e4a778e_u0<=1'h0;
else reg_0e4a778e_u0<=reg_12289738_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00bce4e8_result_delayed_u0<=1'h0;
else reg_00bce4e8_result_delayed_u0<=reg_00bce4e8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_56eb272e_u0<=1'h0;
else reg_56eb272e_u0<=reg_54cc0137_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_710c3541_result_delayed_u0<=1'h0;
else reg_710c3541_result_delayed_u0<=reg_710c3541_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_13e83e22_u0<=1'h0;
else reg_13e83e22_u0<=reg_4ec17b1d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2309bac6_u0<=1'h0;
else reg_2309bac6_u0<=reg_138117ea_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2eae6f7e_u0<=1'h0;
else reg_2eae6f7e_u0<=reg_3b4c4b37_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2e62ff2a_result_delayed_u0<=1'h0;
else reg_2e62ff2a_result_delayed_u0<=reg_2e62ff2a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_63ada2d0_result_delayed_u0<=1'h0;
else reg_63ada2d0_result_delayed_u0<=reg_63ada2d0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_17d8460a_u0<=1'h0;
else reg_17d8460a_u0<=reg_546fd8be_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_63314f9f_result_delayed_u0<=1'h0;
else reg_63314f9f_result_delayed_u0<=reg_63314f9f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_792a283d_result_delayed_u0<=1'h0;
else reg_792a283d_result_delayed_u0<=reg_792a283d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4ec17b1d_u0<=1'h0;
else reg_4ec17b1d_u0<=reg_030c675e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_74e3dda4_result_delayed_u0<=1'h0;
else reg_74e3dda4_result_delayed_u0<=reg_74e3dda4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6cf5c92b_u0<=1'h0;
else reg_6cf5c92b_u0<=reg_6e43fb69_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2cb89c91_result_delayed_u0<=1'h0;
else reg_2cb89c91_result_delayed_u0<=reg_2cb89c91_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1a836fd8_result_delayed_u0<=1'h0;
else reg_1a836fd8_result_delayed_u0<=reg_1a836fd8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3e384fda_u0<=1'h0;
else reg_3e384fda_u0<=reg_01db913f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5fd2d636_u0<=1'h0;
else reg_5fd2d636_u0<=reg_318c1131_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_09c6d144_result_delayed_u0<=1'h0;
else reg_09c6d144_result_delayed_u0<=reg_09c6d144_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_279d2f74_result_delayed_u0<=1'h0;
else reg_279d2f74_result_delayed_u0<=reg_279d2f74_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3b4652ae_u0<=1'h0;
else reg_3b4652ae_u0<=reg_40adac30_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_52747b9c_u0<=1'h0;
else reg_52747b9c_u0<=reg_6f7d9e94_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_689d5d75_u0<=1'h0;
else reg_689d5d75_u0<=reg_7a3ed379_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00bce4e8_result_delayed_result_delayed_u0<=1'h0;
else reg_00bce4e8_result_delayed_result_delayed_u0<=reg_00bce4e8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6f7d9e94_u0<=1'h0;
else reg_6f7d9e94_u0<=reg_37bbd983_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_138117ea_result_delayed_u0<=1'h0;
else reg_138117ea_result_delayed_u0<=reg_138117ea_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5acdfb21_u0<=1'h0;
else reg_5acdfb21_u0<=reg_63daa7a1_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1de599bc_result_delayed_result_delayed_u0<=1'h0;
else reg_1de599bc_result_delayed_result_delayed_u0<=reg_1de599bc_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_030c675e_result_delayed_u0<=1'h0;
else reg_030c675e_result_delayed_u0<=reg_030c675e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_437f3245_result_delayed_u0<=1'h0;
else reg_437f3245_result_delayed_u0<=reg_437f3245_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_63daa7a1_result_delayed_u0<=1'h0;
else reg_63daa7a1_result_delayed_u0<=reg_63daa7a1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_258519cc_result_delayed_result_delayed_u0<=1'h0;
else reg_258519cc_result_delayed_result_delayed_u0<=reg_258519cc_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_158b107d_u0<=1'h0;
else reg_158b107d_u0<=reg_6dc4bd1b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5c74f06b_result_delayed_u0<=1'h0;
else reg_5c74f06b_result_delayed_u0<=reg_5c74f06b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_54cc0137_u0<=1'h0;
else reg_54cc0137_u0<=reg_54826c24_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_57713ae7_result_delayed_u0<=1'h0;
else reg_57713ae7_result_delayed_u0<=reg_57713ae7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0a0626a2_result_delayed_u0<=1'h0;
else reg_0a0626a2_result_delayed_u0<=reg_0a0626a2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_36b55f4a_u0<=1'h0;
else reg_36b55f4a_u0<=reg_6d5cb91c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_05644f67_u0<=1'h0;
else reg_05644f67_u0<=reg_711087ce_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_25493747_u0<=1'h0;
else reg_25493747_u0<=reg_03e66f15_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6741a229_result_delayed_u0<=1'h0;
else reg_6741a229_result_delayed_u0<=reg_6741a229_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_14e9d2f9_u0<=1'h0;
else reg_14e9d2f9_u0<=reg_4e012e31_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7c5e48af_result_delayed_u0<=1'h0;
else reg_7c5e48af_result_delayed_u0<=reg_7c5e48af_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_47eb2b6a_result_delayed_u0<=1'h0;
else reg_47eb2b6a_result_delayed_u0<=reg_47eb2b6a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1de599bc_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_1de599bc_result_delayed_result_delayed_result_delayed_u0<=reg_1de599bc_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7c5e48af_result_delayed_result_delayed_u0<=1'h0;
else reg_7c5e48af_result_delayed_result_delayed_u0<=reg_7c5e48af_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0bd3d5c5_u0<=1'h0;
else reg_0bd3d5c5_u0<=reg_7217fecc_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0e47a050_u0<=1'h0;
else reg_0e47a050_u0<=reg_3b393219_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_76b494ad_u0<=1'h0;
else reg_76b494ad_u0<=reg_515acf62_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_47f4e6ec_result_delayed_u0<=1'h0;
else reg_47f4e6ec_result_delayed_u0<=reg_47f4e6ec_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_792ef732_u0<=1'h0;
else reg_792ef732_u0<=reg_05286558_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_678f3d92_u0<=1'h0;
else reg_678f3d92_u0<=reg_55180568_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_23499f80_result_delayed_u0<=1'h0;
else reg_23499f80_result_delayed_u0<=reg_23499f80_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2309bac6_result_delayed_u0<=1'h0;
else reg_2309bac6_result_delayed_u0<=reg_2309bac6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2ca30e82_u0<=1'h0;
else reg_2ca30e82_u0<=reg_2a1f0d51_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_58bcae9f_u0<=1'h0;
else reg_58bcae9f_u0<=reg_3e784e1c_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_701b11b5_result_delayed_u0<=1'h0;
else reg_701b11b5_result_delayed_u0<=reg_701b11b5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_175ea576_u0<=1'h0;
else reg_175ea576_u0<=reg_062c6117_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0cb5aa9c_u0<=1'h0;
else reg_0cb5aa9c_u0<=reg_13e83e22_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_77dbf5f0_u0<=1'h0;
else reg_77dbf5f0_u0<=reg_6806d06c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5acdfb21_result_delayed_u0<=1'h0;
else reg_5acdfb21_result_delayed_u0<=reg_5acdfb21_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3575e35b_u0<=1'h0;
else reg_3575e35b_u0<=reg_5011c507_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7c5e48af_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_7c5e48af_result_delayed_result_delayed_result_delayed_u0<=reg_7c5e48af_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_18cb5efb_u0<=1'h0;
else reg_18cb5efb_u0<=reg_5f68d729_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_59c65bf7_u0<=1'h0;
else reg_59c65bf7_u0<=reg_41025437_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_701b11b5_result_delayed_result_delayed_u0<=1'h0;
else reg_701b11b5_result_delayed_result_delayed_u0<=reg_701b11b5_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2f53bd66_u0<=1'h0;
else reg_2f53bd66_u0<=reg_3c99258f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4cf96ace_u0<=1'h0;
else reg_4cf96ace_u0<=reg_43039f69_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_33167b6e_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_33167b6e_result_delayed_result_delayed_result_delayed_u0<=reg_33167b6e_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_515acf62_u0<=1'h0;
else reg_515acf62_u0<=reg_44204699_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_37bbd983_u0<=1'h0;
else reg_37bbd983_u0<=reg_682b29b0_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_640558fa_result_delayed_u0<=1'h0;
else reg_640558fa_result_delayed_u0<=reg_640558fa_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7d614f5b_u0<=1'h0;
else reg_7d614f5b_u0<=reg_683a6054_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_78fa2139_result_delayed_u0<=1'h0;
else reg_78fa2139_result_delayed_u0<=reg_78fa2139_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_17699155_u0<=1'h0;
else reg_17699155_u0<=reg_355135b7_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5fd2d636_result_delayed_u0<=1'h0;
else reg_5fd2d636_result_delayed_u0<=reg_5fd2d636_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_09c6d144_result_delayed_result_delayed_u0<=1'h0;
else reg_09c6d144_result_delayed_result_delayed_u0<=reg_09c6d144_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_792a283d_result_delayed_result_delayed_u0<=1'h0;
else reg_792a283d_result_delayed_result_delayed_u0<=reg_792a283d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7dd4b39e_u0<=1'h0;
else reg_7dd4b39e_u0<=reg_78fa2139_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2dac7bf9_u0<=1'h0;
else reg_2dac7bf9_u0<=reg_3c118266_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_107844c4_result_delayed_result_delayed_u0<=1'h0;
else reg_107844c4_result_delayed_result_delayed_u0<=reg_107844c4_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_33b11310_result_delayed_u0<=1'h0;
else reg_33b11310_result_delayed_u0<=reg_33b11310_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5aa7d6c8_result_delayed_u0<=1'h0;
else reg_5aa7d6c8_result_delayed_u0<=reg_5aa7d6c8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_77047715_result_delayed_u0<=1'h0;
else reg_77047715_result_delayed_u0<=reg_77047715_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_03e66f15_result_delayed_u0<=1'h0;
else reg_03e66f15_result_delayed_u0<=reg_03e66f15_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_530b2d69_u0<=1'h0;
else reg_530b2d69_u0<=reg_0c422d83_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0a611af4_result_delayed_u0<=1'h0;
else reg_0a611af4_result_delayed_u0<=reg_0a611af4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3e784e1c_result_delayed_result_delayed_u0<=1'h0;
else reg_3e784e1c_result_delayed_result_delayed_u0<=reg_3e784e1c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5fc6e1a0_u0<=1'h0;
else reg_5fc6e1a0_u0<=reg_32a6867b_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3b393219_result_delayed_u0<=1'h0;
else reg_3b393219_result_delayed_u0<=reg_3b393219_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_70cebea7_u0<=1'h0;
else reg_70cebea7_u0<=reg_5f584dbb_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_31796710_u0<=1'h0;
else reg_31796710_u0<=reg_77dbf5f0_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_370ead64_u0<=1'h0;
else reg_370ead64_u0<=reg_20570b20_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_62f7fc9b_u0<=1'h0;
else reg_62f7fc9b_u0<=reg_297a657a_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_05fe2b93_u0<=1'h0;
else reg_05fe2b93_u0<=reg_536a7781_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01db913f_result_delayed_u0<=1'h0;
else reg_01db913f_result_delayed_u0<=reg_01db913f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3c118266_u0<=1'h0;
else reg_3c118266_u0<=reg_71bdf9cc_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_32fe623a_result_delayed_u0<=1'h0;
else reg_32fe623a_result_delayed_u0<=reg_32fe623a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_387e0416_result_delayed_u0<=1'h0;
else reg_387e0416_result_delayed_u0<=reg_387e0416_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1dd4f50d_result_delayed_u0<=1'h0;
else reg_1dd4f50d_result_delayed_u0<=reg_1dd4f50d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_64870a03_u0<=1'h0;
else reg_64870a03_u0<=reg_1a836fd8_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a88ee59_result_delayed_result_delayed_u0<=1'h0;
else reg_7a88ee59_result_delayed_result_delayed_u0<=reg_7a88ee59_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_485faada_u0<=1'h0;
else reg_485faada_u0<=reg_0a611af4_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7c7216f8_u0<=1'h0;
else reg_7c7216f8_u0<=reg_3d06bf89_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_689528f4_result_delayed_result_delayed_u0<=1'h0;
else reg_689528f4_result_delayed_result_delayed_u0<=reg_689528f4_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u207<=1'h0;
else and_delayed_u207<=and_u3150_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_42afe023_u0<=1'h0;
else reg_42afe023_u0<=reg_4a292b3c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6fbb03a9_result_delayed_result_delayed_u0<=1'h0;
else reg_6fbb03a9_result_delayed_result_delayed_u0<=reg_6fbb03a9_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0a611af4_result_delayed_result_delayed_u0<=1'h0;
else reg_0a611af4_result_delayed_result_delayed_u0<=reg_0a611af4_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_33b11310_result_delayed_result_delayed_u0<=1'h0;
else reg_33b11310_result_delayed_result_delayed_u0<=reg_33b11310_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3d06bf89_u0<=1'h0;
else reg_3d06bf89_u0<=reg_2c3cec3a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_17fed16d_u0<=1'h0;
else reg_17fed16d_u0<=reg_107844c4_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3f347781_result_delayed_u0<=1'h0;
else reg_3f347781_result_delayed_u0<=reg_3f347781_u0;
end
assign mux_u315=(and_u3150_u0)?1'h1:1'h0;
assign or_u895_u0=and_u3150_u0|and_u3149_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_279d2f74_result_delayed_result_delayed_u0<=1'h0;
else reg_279d2f74_result_delayed_result_delayed_u0<=reg_279d2f74_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_54cc0137_result_delayed_u0<=1'h0;
else reg_54cc0137_result_delayed_u0<=reg_54cc0137_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_27e96f4d_result_delayed_result_delayed_u0<=1'h0;
else reg_27e96f4d_result_delayed_result_delayed_u0<=reg_27e96f4d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_57b67e1e_result_delayed_u0<=1'h0;
else reg_57b67e1e_result_delayed_u0<=reg_57b67e1e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_355135b7_result_delayed_result_delayed_u0<=1'h0;
else reg_355135b7_result_delayed_result_delayed_u0<=reg_355135b7_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1536340b_result_delayed_u0<=1'h0;
else reg_1536340b_result_delayed_u0<=reg_1536340b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3c99258f_result_delayed_u0<=1'h0;
else reg_3c99258f_result_delayed_u0<=reg_3c99258f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_05fe2b93_result_delayed_u0<=1'h0;
else reg_05fe2b93_result_delayed_u0<=reg_05fe2b93_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4b516dfb_u0<=1'h0;
else reg_4b516dfb_u0<=reg_0a6e669d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6e43fb69_result_delayed_u0<=1'h0;
else reg_6e43fb69_result_delayed_u0<=reg_6e43fb69_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7c7f1881_result_delayed_u0<=1'h0;
else reg_7c7f1881_result_delayed_u0<=reg_7c7f1881_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_04854db4_result_delayed_u0<=1'h0;
else reg_04854db4_result_delayed_u0<=reg_04854db4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3e384fda_result_delayed_u0<=1'h0;
else reg_3e384fda_result_delayed_u0<=reg_3e384fda_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_09c6d144_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_09c6d144_result_delayed_result_delayed_result_delayed_u0<=reg_09c6d144_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3715a5a1_u0<=1'h0;
else reg_3715a5a1_u0<=reg_0304da20_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_33b11310_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_33b11310_result_delayed_result_delayed_result_delayed_u0<=reg_33b11310_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_62f7fc9b_result_delayed_u0<=1'h0;
else reg_62f7fc9b_result_delayed_u0<=reg_62f7fc9b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_54fa2642_u0<=1'h0;
else reg_54fa2642_u0<=reg_32e22ff9_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_44204699_u0<=1'h0;
else reg_44204699_u0<=reg_7bc1bfcd_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_03ce3977_u0<=1'h0;
else reg_03ce3977_u0<=reg_40e76b7d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_28399a83_u0<=1'h0;
else reg_28399a83_u0<=reg_05fa154c_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_57713ae7_result_delayed_result_delayed_u0<=1'h0;
else reg_57713ae7_result_delayed_result_delayed_u0<=reg_57713ae7_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2ecaeed5_result_delayed_result_delayed_u0<=1'h0;
else reg_2ecaeed5_result_delayed_result_delayed_u0<=reg_2ecaeed5_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2a1c2b8c_result_delayed_u0<=1'h0;
else reg_2a1c2b8c_result_delayed_u0<=reg_2a1c2b8c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_78fa2139_result_delayed_result_delayed_u0<=1'h0;
else reg_78fa2139_result_delayed_result_delayed_u0<=reg_78fa2139_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a88ee59_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_7a88ee59_result_delayed_result_delayed_result_delayed_u0<=reg_7a88ee59_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_40adac30_result_delayed_result_delayed_u0<=1'h0;
else reg_40adac30_result_delayed_result_delayed_u0<=reg_40adac30_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2dac7bf9_result_delayed_u0<=1'h0;
else reg_2dac7bf9_result_delayed_u0<=reg_2dac7bf9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5085924e_u0<=1'h0;
else reg_5085924e_u0<=reg_770cdc1d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6d657fae_u0<=1'h0;
else reg_6d657fae_u0<=reg_7b23ef69_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_05074d01_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_05074d01_result_delayed_result_delayed_result_delayed_u0<=reg_05074d01_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_18cb5efb_result_delayed_u0<=1'h0;
else reg_18cb5efb_result_delayed_u0<=reg_18cb5efb_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_77b9b56b_u0<=1'h0;
else reg_77b9b56b_u0<=reg_1536340b_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7bc1bfcd_result_delayed_u0<=1'h0;
else reg_7bc1bfcd_result_delayed_u0<=reg_7bc1bfcd_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0edfde7a_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_0edfde7a_result_delayed_result_delayed_result_delayed_u0<=reg_0edfde7a_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2c3cec3a_result_delayed_u0<=1'h0;
else reg_2c3cec3a_result_delayed_u0<=reg_2c3cec3a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5fc6e1a0_result_delayed_u0<=1'h0;
else reg_5fc6e1a0_result_delayed_u0<=reg_5fc6e1a0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_107844c4_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_107844c4_result_delayed_result_delayed_result_delayed_u0<=reg_107844c4_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2349ca1b_result_delayed_u0<=1'h0;
else reg_2349ca1b_result_delayed_u0<=reg_2349ca1b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4d6a0c19_result_delayed_u0<=1'h0;
else reg_4d6a0c19_result_delayed_u0<=reg_4d6a0c19_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_546fd8be_result_delayed_u0<=1'h0;
else reg_546fd8be_result_delayed_u0<=reg_546fd8be_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2c075897_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_2c075897_result_delayed_result_delayed_result_delayed_u0<=reg_2c075897_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_57b67e1e_result_delayed_result_delayed_u0<=1'h0;
else reg_57b67e1e_result_delayed_result_delayed_u0<=reg_57b67e1e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_429ea278_result_delayed_u0<=1'h0;
else reg_429ea278_result_delayed_u0<=reg_429ea278_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_711087ce_u0<=1'h0;
else reg_711087ce_u0<=reg_3715a5a1_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2d3a4979_result_delayed_u0<=1'h0;
else reg_2d3a4979_result_delayed_u0<=reg_2d3a4979_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5f584dbb_u0<=1'h0;
else reg_5f584dbb_u0<=reg_049d2474_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_35da391c_result_delayed_u0<=1'h0;
else reg_35da391c_result_delayed_u0<=reg_35da391c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_258519cc_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_258519cc_result_delayed_result_delayed_result_delayed_u0<=reg_258519cc_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_13e83e22_result_delayed_u0<=1'h0;
else reg_13e83e22_result_delayed_u0<=reg_13e83e22_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_43b7c159_u0<=1'h0;
else reg_43b7c159_u0<=reg_5780a32a_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00326d3c_result_delayed_result_delayed_u0<=1'h0;
else reg_00326d3c_result_delayed_result_delayed_u0<=reg_00326d3c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1de599bc_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_1de599bc_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_1de599bc_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_71bdf9cc_result_delayed_u0<=1'h0;
else reg_71bdf9cc_result_delayed_u0<=reg_71bdf9cc_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1a836fd8_result_delayed_result_delayed_u0<=1'h0;
else reg_1a836fd8_result_delayed_result_delayed_u0<=reg_1a836fd8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2ca30e82_result_delayed_u0<=1'h0;
else reg_2ca30e82_result_delayed_u0<=reg_2ca30e82_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5b15db0b_result_delayed_u0<=1'h0;
else reg_5b15db0b_result_delayed_u0<=reg_5b15db0b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0a6e669d_result_delayed_u0<=1'h0;
else reg_0a6e669d_result_delayed_u0<=reg_0a6e669d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_54cc0137_result_delayed_result_delayed_u0<=1'h0;
else reg_54cc0137_result_delayed_result_delayed_u0<=reg_54cc0137_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2eae6f7e_result_delayed_u0<=1'h0;
else reg_2eae6f7e_result_delayed_u0<=reg_2eae6f7e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0fb3eac1_result_delayed_u0<=1'h0;
else reg_0fb3eac1_result_delayed_u0<=reg_0fb3eac1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5011c507_result_delayed_u0<=1'h0;
else reg_5011c507_result_delayed_u0<=reg_5011c507_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_32e22ff9_result_delayed_u0<=1'h0;
else reg_32e22ff9_result_delayed_u0<=reg_32e22ff9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_43d5e336_result_delayed_u0<=1'h0;
else reg_43d5e336_result_delayed_u0<=reg_43d5e336_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_05286558_result_delayed_u0<=1'h0;
else reg_05286558_result_delayed_u0<=reg_05286558_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_14e9d2f9_result_delayed_u0<=1'h0;
else reg_14e9d2f9_result_delayed_u0<=reg_14e9d2f9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5d8c3e8b_u0<=1'h0;
else reg_5d8c3e8b_u0<=reg_33b11310_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0bfe7f33_result_delayed_u0<=1'h0;
else reg_0bfe7f33_result_delayed_u0<=reg_0bfe7f33_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_05fe2b93_result_delayed_result_delayed_u0<=1'h0;
else reg_05fe2b93_result_delayed_result_delayed_u0<=reg_05fe2b93_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_03e66f15_result_delayed_result_delayed_u0<=1'h0;
else reg_03e66f15_result_delayed_result_delayed_u0<=reg_03e66f15_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_50917495_result_delayed_u0<=1'h0;
else reg_50917495_result_delayed_u0<=reg_50917495_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_770cdc1d_u0<=1'h0;
else reg_770cdc1d_u0<=reg_7a51229e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_258519cc_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_258519cc_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_258519cc_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7b23ef69_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_7b23ef69_result_delayed_result_delayed_result_delayed_u0<=reg_7b23ef69_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_09c6d144_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_09c6d144_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_09c6d144_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5c72dd07_result_delayed_u0<=1'h0;
else reg_5c72dd07_result_delayed_u0<=reg_5c72dd07_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_77dbf5f0_result_delayed_u0<=1'h0;
else reg_77dbf5f0_result_delayed_u0<=reg_77dbf5f0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1536340b_result_delayed_result_delayed_u0<=1'h0;
else reg_1536340b_result_delayed_result_delayed_u0<=reg_1536340b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0304da20_result_delayed_result_delayed_u0<=1'h0;
else reg_0304da20_result_delayed_result_delayed_u0<=reg_0304da20_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_401b0405_result_delayed_u0<=1'h0;
else reg_401b0405_result_delayed_u0<=reg_401b0405_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_50917495_result_delayed_result_delayed_u0<=1'h0;
else reg_50917495_result_delayed_result_delayed_u0<=reg_50917495_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_682b29b0_result_delayed_u0<=1'h0;
else reg_682b29b0_result_delayed_u0<=reg_682b29b0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a3ed379_result_delayed_u0<=1'h0;
else reg_7a3ed379_result_delayed_u0<=reg_7a3ed379_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_66095291_result_delayed_u0<=1'h0;
else reg_66095291_result_delayed_u0<=reg_66095291_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7ec4fde8_u0<=1'h0;
else reg_7ec4fde8_u0<=reg_1ca67dbd_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0e12093d_u0<=1'h0;
else reg_0e12093d_u0<=reg_3d4ff93c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_689528f4_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_689528f4_result_delayed_result_delayed_result_delayed_u0<=reg_689528f4_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0c422d83_result_delayed_u0<=1'h0;
else reg_0c422d83_result_delayed_u0<=reg_0c422d83_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_31796710_result_delayed_u0<=1'h0;
else reg_31796710_result_delayed_u0<=reg_31796710_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_062c6117_u0<=1'h0;
else reg_062c6117_u0<=reg_7ec4fde8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_41025437_result_delayed_u0<=1'h0;
else reg_41025437_result_delayed_u0<=reg_41025437_u0;
end
assign and_u3151_u0=and_u3146_u0&and_u3152_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5fd2d636_result_delayed_result_delayed_u0<=1'h0;
else reg_5fd2d636_result_delayed_result_delayed_u0<=reg_5fd2d636_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_23b56b6a_result_delayed_u0<=1'h0;
else reg_23b56b6a_result_delayed_u0<=reg_23b56b6a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_318c1131_result_delayed_u0<=1'h0;
else reg_318c1131_result_delayed_u0<=reg_318c1131_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_638aaf04_result_delayed_u0<=1'h0;
else reg_638aaf04_result_delayed_u0<=reg_638aaf04_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_74c8f38e_u0<=1'h0;
else reg_74c8f38e_u0<=reg_77b9b56b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_638aaf04_result_delayed_result_delayed_u0<=1'h0;
else reg_638aaf04_result_delayed_result_delayed_u0<=reg_638aaf04_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_41bcb2f2_u0<=1'h0;
else reg_41bcb2f2_u0<=reg_64fa00de_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2a1f0d51_u0<=1'h0;
else reg_2a1f0d51_u0<=reg_0bfe7f33_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1ca67dbd_result_delayed_u0<=1'h0;
else reg_1ca67dbd_result_delayed_u0<=reg_1ca67dbd_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_63daa7a1_result_delayed_result_delayed_u0<=1'h0;
else reg_63daa7a1_result_delayed_result_delayed_u0<=reg_63daa7a1_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_05fa154c_result_delayed_result_delayed_u0<=1'h0;
else reg_05fa154c_result_delayed_result_delayed_u0<=reg_05fa154c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_37bbd983_result_delayed_u0<=1'h0;
else reg_37bbd983_result_delayed_u0<=reg_37bbd983_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6741a229_result_delayed_result_delayed_u0<=1'h0;
else reg_6741a229_result_delayed_result_delayed_u0<=reg_6741a229_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6741a229_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_6741a229_result_delayed_result_delayed_result_delayed_u0<=reg_6741a229_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1db07eea_u0<=1'h0;
else reg_1db07eea_u0<=reg_7f7d622f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0afd59a6_u0<=1'h0;
else reg_0afd59a6_u0<=reg_792a283d_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0e12093d_result_delayed_u0<=1'h0;
else reg_0e12093d_result_delayed_u0<=reg_0e12093d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_15387666_u0<=1'h0;
else reg_15387666_u0<=reg_29782e98_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5780a32a_result_delayed_u0<=1'h0;
else reg_5780a32a_result_delayed_u0<=reg_5780a32a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3ac681a6_u0<=1'h0;
else reg_3ac681a6_u0<=reg_1536c80b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_792a283d_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_792a283d_result_delayed_result_delayed_result_delayed_u0<=reg_792a283d_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_64870a03_result_delayed_u0<=1'h0;
else reg_64870a03_result_delayed_u0<=reg_64870a03_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_678f3d92_result_delayed_u0<=1'h0;
else reg_678f3d92_result_delayed_u0<=reg_678f3d92_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_387e0416_result_delayed_result_delayed_u0<=1'h0;
else reg_387e0416_result_delayed_result_delayed_u0<=reg_387e0416_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_049d2474_result_delayed_u0<=1'h0;
else reg_049d2474_result_delayed_u0<=reg_049d2474_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_711087ce_result_delayed_u0<=1'h0;
else reg_711087ce_result_delayed_u0<=reg_711087ce_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3b4c4b37_result_delayed_u0<=1'h0;
else reg_3b4c4b37_result_delayed_u0<=reg_3b4c4b37_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_33b11310_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_33b11310_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_33b11310_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_20570b20_u0<=1'h0;
else reg_20570b20_u0<=reg_17e75387_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_37bbd983_result_delayed_result_delayed_u0<=1'h0;
else reg_37bbd983_result_delayed_result_delayed_u0<=reg_37bbd983_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2a1f0d51_result_delayed_u0<=1'h0;
else reg_2a1f0d51_result_delayed_u0<=reg_2a1f0d51_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_55180568_result_delayed_u0<=1'h0;
else reg_55180568_result_delayed_u0<=reg_55180568_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_70cebea7_result_delayed_u0<=1'h0;
else reg_70cebea7_result_delayed_u0<=reg_70cebea7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_297a657a_result_delayed_u0<=1'h0;
else reg_297a657a_result_delayed_u0<=reg_297a657a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5aa7d6c8_result_delayed_result_delayed_u0<=1'h0;
else reg_5aa7d6c8_result_delayed_result_delayed_u0<=reg_5aa7d6c8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_47f4e6ec_result_delayed_result_delayed_u0<=1'h0;
else reg_47f4e6ec_result_delayed_result_delayed_u0<=reg_47f4e6ec_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1b8047bd_result_delayed_u0<=1'h0;
else reg_1b8047bd_result_delayed_u0<=reg_1b8047bd_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7f7d622f_result_delayed_u0<=1'h0;
else reg_7f7d622f_result_delayed_u0<=reg_7f7d622f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5011c507_result_delayed_result_delayed_u0<=1'h0;
else reg_5011c507_result_delayed_result_delayed_u0<=reg_5011c507_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_539db809_u0<=1'h0;
else reg_539db809_u0<=reg_6109ede1_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0bfe7f33_result_delayed_result_delayed_u0<=1'h0;
else reg_0bfe7f33_result_delayed_result_delayed_u0<=reg_0bfe7f33_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_40e76b7d_u0<=1'h0;
else reg_40e76b7d_u0<=reg_7ff55f76_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_40d160ea_result_delayed_u0<=1'h0;
else reg_40d160ea_result_delayed_u0<=reg_40d160ea_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7217fecc_result_delayed_u0<=1'h0;
else reg_7217fecc_result_delayed_u0<=reg_7217fecc_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4e012e31_result_delayed_u0<=1'h0;
else reg_4e012e31_result_delayed_u0<=reg_4e012e31_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7ff55f76_result_delayed_result_delayed_u0<=1'h0;
else reg_7ff55f76_result_delayed_result_delayed_u0<=reg_7ff55f76_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6d5cb91c_result_delayed_u0<=1'h0;
else reg_6d5cb91c_result_delayed_u0<=reg_6d5cb91c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5f68d729_result_delayed_u0<=1'h0;
else reg_5f68d729_result_delayed_u0<=reg_5f68d729_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3715a5a1_result_delayed_u0<=1'h0;
else reg_3715a5a1_result_delayed_u0<=reg_3715a5a1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_41025437_result_delayed_result_delayed_u0<=1'h0;
else reg_41025437_result_delayed_result_delayed_u0<=reg_41025437_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6109ede1_result_delayed_u0<=1'h0;
else reg_6109ede1_result_delayed_u0<=reg_6109ede1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4a292b3c_result_delayed_u0<=1'h0;
else reg_4a292b3c_result_delayed_u0<=reg_4a292b3c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7ec4fde8_result_delayed_u0<=1'h0;
else reg_7ec4fde8_result_delayed_u0<=reg_7ec4fde8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_378e778c_result_delayed_u0<=1'h0;
else reg_378e778c_result_delayed_u0<=reg_378e778c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_64fa00de_result_delayed_result_delayed_u0<=1'h0;
else reg_64fa00de_result_delayed_result_delayed_u0<=reg_64fa00de_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0e47a050_result_delayed_u0<=1'h0;
else reg_0e47a050_result_delayed_u0<=reg_0e47a050_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_17e75387_result_delayed_u0<=1'h0;
else reg_17e75387_result_delayed_u0<=reg_17e75387_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3d4ff93c_result_delayed_u0<=1'h0;
else reg_3d4ff93c_result_delayed_u0<=reg_3d4ff93c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_15387666_result_delayed_u0<=1'h0;
else reg_15387666_result_delayed_u0<=reg_15387666_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_12289738_result_delayed_u0<=1'h0;
else reg_12289738_result_delayed_u0<=reg_12289738_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_74e3dda4_result_delayed_result_delayed_u0<=1'h0;
else reg_74e3dda4_result_delayed_result_delayed_u0<=reg_74e3dda4_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4b39e741_result_delayed_u0<=1'h0;
else reg_4b39e741_result_delayed_u0<=reg_4b39e741_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_54826c24_result_delayed_u0<=1'h0;
else reg_54826c24_result_delayed_u0<=reg_54826c24_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_297a657a_result_delayed_result_delayed_u0<=1'h0;
else reg_297a657a_result_delayed_result_delayed_u0<=reg_297a657a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6806d06c_result_delayed_u0<=1'h0;
else reg_6806d06c_result_delayed_u0<=reg_6806d06c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0c3478e6_result_delayed_result_delayed_u0<=1'h0;
else reg_0c3478e6_result_delayed_result_delayed_u0<=reg_0c3478e6_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1536c80b_result_delayed_u0<=1'h0;
else reg_1536c80b_result_delayed_u0<=reg_1536c80b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a51229e_result_delayed_u0<=1'h0;
else reg_7a51229e_result_delayed_u0<=reg_7a51229e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6dc4bd1b_result_delayed_u0<=1'h0;
else reg_6dc4bd1b_result_delayed_u0<=reg_6dc4bd1b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_43039f69_result_delayed_result_delayed_u0<=1'h0;
else reg_43039f69_result_delayed_result_delayed_u0<=reg_43039f69_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5780a32a_result_delayed_result_delayed_u0<=1'h0;
else reg_5780a32a_result_delayed_result_delayed_u0<=reg_5780a32a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_29782e98_u0<=1'h0;
else reg_29782e98_u0<=reg_35ff7cc6_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_536a7781_result_delayed_u0<=1'h0;
else reg_536a7781_result_delayed_u0<=reg_536a7781_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_32a6867b_result_delayed_result_delayed_u0<=1'h0;
else reg_32a6867b_result_delayed_result_delayed_u0<=reg_32a6867b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_683a6054_result_delayed_u0<=1'h0;
else reg_683a6054_result_delayed_u0<=reg_683a6054_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_58bcae9f_result_delayed_u0<=1'h0;
else reg_58bcae9f_result_delayed_u0<=reg_58bcae9f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7d614f5b_result_delayed_u0<=1'h0;
else reg_7d614f5b_result_delayed_u0<=reg_7d614f5b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_57b67e1e_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_57b67e1e_result_delayed_result_delayed_result_delayed_u0<=reg_57b67e1e_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4cf96ace_result_delayed_u0<=1'h0;
else reg_4cf96ace_result_delayed_u0<=reg_4cf96ace_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_35ff7cc6_result_delayed_u0<=1'h0;
else reg_35ff7cc6_result_delayed_u0<=reg_35ff7cc6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u208_u0<=1'h0;
else and_delayed_u208_u0<=and_u3151_u0;
end
assign or_u896_u0=reg_23499f80_result_delayed_u0|and_delayed_u208_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_77b9b56b_result_delayed_u0<=1'h0;
else reg_77b9b56b_result_delayed_u0<=reg_77b9b56b_u0;
end
assign or_u897_u0=and_u3153_u0|and_u3150_u0;
assign and_u3152_u0=and_u3143_u0&and_u3155_u0;
assign and_u3153_u0=and_u3144_u0&and_u3155_u0;
assign or_u898_u0=and_u3153_u0|or_u895_u0;
assign mux_u316_u0=(and_u3153_u0)?1'h1:mux_u315;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_58165587_u0<=1'h0;
else reg_58165587_u0<=reg_31cf41da_u0;
end
assign or_u899_u0=and_u3153_u0|and_u3150_u0;
assign mux_u317_u0=(and_u3153_u0)?32'h2:32'h200;
assign or_u900_u0=and_u3153_u0|and_u3150_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_31cf41da_u0<=1'h0;
else reg_31cf41da_u0<=and_delayed_u209_u0;
end
assign or_u901_u0=and_u3153_u0|and_u3150_u0;
assign or_u902_u0=reg_58165587_u0|or_u896_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u209_u0<=1'h0;
else and_delayed_u209_u0<=and_u3153_u0;
end
assign and_u3154_u0=and_u3141_u0&and_u3140_u0;
assign and_u3155_u0=and_u3142_u0&and_u3140_u0;
assign or_u903_u0=or_u902_u0|and_delayed_u210_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u210_u0<=1'h0;
else and_delayed_u210_u0<=and_u3154_u0;
end
assign equals_u166_a_signed={31'b0, port_0a81f2c6_};
assign equals_u166_b_signed=32'h1;
assign equals_u166=equals_u166_a_signed==equals_u166_b_signed;
assign and_u3156_u0=and_u3140_u0&equals_u166;
assign not_u530_u0=~equals_u166;
assign and_u3157_u0=and_u3140_u0&not_u530_u0;
assign and_u3158_u0=and_u3172_u0&port_5071c1a7_;
assign not_u531_u0=~port_5071c1a7_;
assign and_u3159_u0=and_u3172_u0&not_u531_u0;
assign lessThan_u75_a_signed=port_3bb784d0_;
assign lessThan_u75_b_signed=port_1ca215c6_;
assign lessThan_u75=lessThan_u75_a_signed<lessThan_u75_b_signed;
assign and_u3160_u0=and_u3169_u0&lessThan_u75;
assign and_u3161_u0=and_u3169_u0&not_u532_u0;
assign not_u532_u0=~lessThan_u75;
assign and_u3162_u0=and_u3168_u0&port_2adbeb14_;
assign and_u3163_u0=and_u3168_u0&not_u533_u0;
assign not_u533_u0=~port_2adbeb14_;
assign add=port_3bb784d0_+32'h0;
assign and_u3164_u0=and_u3166_u0&port_63d562ec_;
assign simplePinWrite_u468=16'h1&{16{1'h1}};
assign simplePinWrite_u469=port_2ccab656_;
assign simplePinWrite_u470=and_u3166_u0&{1{and_u3166_u0}};
assign add_u374=port_3bb784d0_+32'h1;
always @(posedge CLK)
begin
if (and_u3166_u0)
syncEnable_u550<=port_2ccab656_;
end
assign and_u3165_u0=and_u3163_u0&and_u3168_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0de2a3c0_u0<=1'h0;
else reg_0de2a3c0_u0<=and_u3166_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u211_u0<=1'h0;
else and_delayed_u211_u0<=and_u3165_u0;
end
assign mux_u318_u0=(reg_0de2a3c0_u0)?syncEnable_u550:syncEnable_u551_u0;
always @(posedge CLK)
begin
if (and_u3168_u0)
syncEnable_u551_u0<=mux_u329_u0;
end
assign and_u3166_u0=and_u3162_u0&and_u3168_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0498419c_u0<=1'h0;
else reg_0498419c_u0<=and_u3168_u0;
end
assign mux_u319_u0=(reg_0498419c_u0)?mux_u318_u0:syncEnable_u553_u0;
assign mux_u320_u0=(reg_0498419c_u0)?syncEnable_u552_u0:32'h0;
always @(posedge CLK)
begin
if (and_u3169_u0)
syncEnable_u552_u0<=mux_u330_u0;
end
always @(posedge CLK)
begin
if (and_u3169_u0)
syncEnable_u553_u0<=mux_u329_u0;
end
assign and_u3167_u0=and_u3161_u0&and_u3169_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u212_u0<=1'h0;
else and_delayed_u212_u0<=and_u3167_u0;
end
assign and_u3168_u0=and_u3160_u0&and_u3169_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_490a59eb_u0<=1'h0;
else reg_490a59eb_u0<=and_u3170_u0;
end
assign mux_u321_u0=(reg_490a59eb_u0)?syncEnable_u554_u0:mux_u319_u0;
assign mux_u322_u0=(reg_490a59eb_u0)?syncEnable_u555_u0:mux_u320_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5602ca0c_u0<=1'h0;
else reg_5602ca0c_u0<=and_u3169_u0;
end
assign and_u3169_u0=and_u3158_u0&and_u3172_u0;
always @(posedge CLK)
begin
if (and_u3172_u0)
syncEnable_u554_u0<=mux_u329_u0;
end
always @(posedge CLK)
begin
if (and_u3172_u0)
syncEnable_u555_u0<=mux_u330_u0;
end
assign and_u3170_u0=and_u3159_u0&and_u3172_u0;
assign mux_u323_u0=(and_delayed_u213_u0)?syncEnable_u557_u0:mux_u321_u0;
assign and_u3171_u0=and_u3157_u0&and_u3140_u0;
always @(posedge CLK)
begin
if (and_u3140_u0)
syncEnable_u556_u0<=mux_u330_u0;
end
assign mux_u324_u0=(and_delayed_u213_u0)?syncEnable_u556_u0:mux_u322_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7e9a4e4d_u0<=1'h0;
else reg_7e9a4e4d_u0<=and_u3172_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u213_u0<=1'h0;
else and_delayed_u213_u0<=and_u3171_u0;
end
assign and_u3172_u0=and_u3156_u0&and_u3140_u0;
always @(posedge CLK)
begin
if (and_u3140_u0)
syncEnable_u557_u0<=mux_u329_u0;
end
always @(posedge CLK)
begin
if (block_GO_delayed_u10)
latch_3dab8262_reg<=mux_u323_u0;
end
assign latch_3dab8262_out=(block_GO_delayed_u10)?mux_u323_u0:latch_3dab8262_reg;
assign mux_u325_u0=(or_u899_u0)?1'h1:1'h0;
assign or_u904_u0=or_u899_u0|and_u3167_u0;
assign or_u905_u0=or_u898_u0|and_u3167_u0;
assign mux_u326_u0=(or_u898_u0)?mux_u316_u0:1'h0;
always @(posedge CLK)
begin
if (block_GO_delayed_u10)
latch_182feb1c_reg<=mux_u324_u0;
end
assign latch_182feb1c_out=(block_GO_delayed_u10)?mux_u324_u0:latch_182feb1c_reg;
assign mux_u327_u0=(or_u900_u0)?{22'b0, mux_u317_u0[9], 7'b0, mux_u317_u0[1], 1'b0}:32'hffffffff;
assign or_u906_u0=or_u900_u0|and_u3167_u0;
assign mux_u328_u0=(or_u897_u0)?32'h0:add_u374;
assign or_u907_u0=or_u897_u0|and_u3166_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
block_GO_delayed_u10<=1'h0;
else block_GO_delayed_u10<=and_u3140_u0;
end
always @(posedge CLK)
begin
if (or_u903_u0)
fbReg_temp_fsmOldState_resized_LH1_xy_6_u0<=latch_182feb1c_out;
end
assign mux_u329_u0=(reg_687233e3_result_delayed_u0)?16'h0:fbReg_Out1Portvalue_u3;
assign mux_u330_u0=(reg_687233e3_result_delayed_u0)?32'h0:fbReg_temp_fsmOldState_resized_LH1_xy_6_u0;
always @(posedge CLK)
begin
if (or_u903_u0)
fbReg_Out1Portvalue_u3<=latch_3dab8262_out;
end
always @(posedge CLK)
begin
if (reg_687233e3_result_delayed_u0)
syncEnable_u558_u0<=RESET;
end
always @(posedge CLK or posedge syncEnable_u558_u0)
begin
if (syncEnable_u558_u0)
loopControl_u7<=1'h0;
else loopControl_u7<=or_u903_u0;
end
assign or_u908_u0=reg_687233e3_result_delayed_u0|loopControl_u7;
assign mux_u331_u0=(GO)?32'h0:mux_u328_u0;
assign or_u909_u0=GO|or_u907_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_687233e3_u0<=1'h0;
else reg_687233e3_u0<=GO;
end
assign or_u910_u0=GO|or_u901_u0;
assign mux_u332_u0=(GO)?1'h0:mux_u326_u0;
assign or_u911_u0=GO|or_u905_u0;
assign mux_u333_u0=(GO)?1'h0:mux_u325_u0;
assign or_u912_u0=GO|or_u904_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_687233e3_result_delayed_u0<=1'h0;
else reg_687233e3_result_delayed_u0<=reg_687233e3_u0;
end
assign mux_u334_u0=(GO)?32'hffffffff:mux_u327_u0;
assign or_u913_u0=GO|or_u906_u0;
assign RESULT=or_u910_u0;
assign RESULT_u1863=32'h0;
assign RESULT_u1864=or_u911_u0;
assign RESULT_u1865=mux_u332_u0;
assign RESULT_u1866=or_u909_u0;
assign RESULT_u1867=mux_u331_u0;
assign RESULT_u1868=or_u913_u0;
assign RESULT_u1869=mux_u334_u0;
assign RESULT_u1870=or_u912_u0;
assign RESULT_u1871=mux_u333_u0;
assign RESULT_u1872=and_u3166_u0;
assign RESULT_u1873=add;
assign RESULT_u1874=3'h1;
assign RESULT_u1875=simplePinWrite;
assign RESULT_u1876=simplePinWrite_u468;
assign RESULT_u1877=simplePinWrite_u466;
assign RESULT_u1878=simplePinWrite_u467;
assign RESULT_u1879=simplePinWrite_u469;
assign RESULT_u1880=simplePinWrite_u470;
assign DONE=1'h0;
endmodule



module resized_LH1_xy_endianswapper_0a8130a3_(endianswapper_0a8130a3_in, endianswapper_0a8130a3_out);
input	[31:0]	endianswapper_0a8130a3_in;
output	[31:0]	endianswapper_0a8130a3_out;
assign endianswapper_0a8130a3_out=endianswapper_0a8130a3_in;
endmodule



module resized_LH1_xy_endianswapper_222b5ae4_(endianswapper_222b5ae4_in, endianswapper_222b5ae4_out);
input	[31:0]	endianswapper_222b5ae4_in;
output	[31:0]	endianswapper_222b5ae4_out;
assign endianswapper_222b5ae4_out=endianswapper_222b5ae4_in;
endmodule



module resized_LH1_xy_stateVar_Out1TokenIndex(bus_44763466_, bus_08eb61b0_, bus_3d7dc20a_, bus_1be81a8d_, bus_4a96edb8_);
input		bus_44763466_;
input		bus_08eb61b0_;
input		bus_3d7dc20a_;
input	[31:0]	bus_1be81a8d_;
output	[31:0]	bus_4a96edb8_;
reg	[31:0]	stateVar_Out1TokenIndex_u3=32'h0;
wire	[31:0]	endianswapper_0a8130a3_out;
wire	[31:0]	endianswapper_222b5ae4_out;
always @(posedge bus_44763466_ or posedge bus_08eb61b0_)
begin
if (bus_08eb61b0_)
stateVar_Out1TokenIndex_u3<=32'h0;
else if (bus_3d7dc20a_)
stateVar_Out1TokenIndex_u3<=endianswapper_0a8130a3_out;
end
resized_LH1_xy_endianswapper_0a8130a3_ resized_LH1_xy_endianswapper_0a8130a3__1(.endianswapper_0a8130a3_in(bus_1be81a8d_), 
  .endianswapper_0a8130a3_out(endianswapper_0a8130a3_out));
assign bus_4a96edb8_=endianswapper_222b5ae4_out;
resized_LH1_xy_endianswapper_222b5ae4_ resized_LH1_xy_endianswapper_222b5ae4__1(.endianswapper_222b5ae4_in(stateVar_Out1TokenIndex_u3), 
  .endianswapper_222b5ae4_out(endianswapper_222b5ae4_out));
endmodule



module resized_LH1_xy_endianswapper_2275df71_(endianswapper_2275df71_in, endianswapper_2275df71_out);
input	[31:0]	endianswapper_2275df71_in;
output	[31:0]	endianswapper_2275df71_out;
assign endianswapper_2275df71_out=endianswapper_2275df71_in;
endmodule



module resized_LH1_xy_endianswapper_7eb888e7_(endianswapper_7eb888e7_in, endianswapper_7eb888e7_out);
input	[31:0]	endianswapper_7eb888e7_in;
output	[31:0]	endianswapper_7eb888e7_out;
assign endianswapper_7eb888e7_out=endianswapper_7eb888e7_in;
endmodule



module resized_LH1_xy_stateVar_Out1MaxTokenIndex(bus_344cf808_, bus_2e472a30_, bus_463825f8_, bus_02e6a7a9_, bus_7668b64d_);
input		bus_344cf808_;
input		bus_2e472a30_;
input		bus_463825f8_;
input	[31:0]	bus_02e6a7a9_;
output	[31:0]	bus_7668b64d_;
wire	[31:0]	endianswapper_2275df71_out;
reg	[31:0]	stateVar_Out1MaxTokenIndex_u3=32'h0;
wire	[31:0]	endianswapper_7eb888e7_out;
resized_LH1_xy_endianswapper_2275df71_ resized_LH1_xy_endianswapper_2275df71__1(.endianswapper_2275df71_in(bus_02e6a7a9_), 
  .endianswapper_2275df71_out(endianswapper_2275df71_out));
assign bus_7668b64d_=endianswapper_7eb888e7_out;
always @(posedge bus_344cf808_ or posedge bus_2e472a30_)
begin
if (bus_2e472a30_)
stateVar_Out1MaxTokenIndex_u3<=32'h0;
else if (bus_463825f8_)
stateVar_Out1MaxTokenIndex_u3<=endianswapper_2275df71_out;
end
resized_LH1_xy_endianswapper_7eb888e7_ resized_LH1_xy_endianswapper_7eb888e7__1(.endianswapper_7eb888e7_in(stateVar_Out1MaxTokenIndex_u3), 
  .endianswapper_7eb888e7_out(endianswapper_7eb888e7_out));
endmodule



module resized_LH1_xy_endianswapper_6acb6654_(endianswapper_6acb6654_in, endianswapper_6acb6654_out);
input	[15:0]	endianswapper_6acb6654_in;
output	[15:0]	endianswapper_6acb6654_out;
assign endianswapper_6acb6654_out=endianswapper_6acb6654_in;
endmodule



module resized_LH1_xy_endianswapper_34cf1120_(endianswapper_34cf1120_in, endianswapper_34cf1120_out);
input	[15:0]	endianswapper_34cf1120_in;
output	[15:0]	endianswapper_34cf1120_out;
assign endianswapper_34cf1120_out=endianswapper_34cf1120_in;
endmodule



module resized_LH1_xy_stateVar_rowRepeated(bus_1d013d35_, bus_1beb5227_, bus_0469fc4f_, bus_51ae933d_, bus_6a8dff02_, bus_733d2b23_, bus_70ada90a_);
input		bus_1d013d35_;
input		bus_1beb5227_;
input		bus_0469fc4f_;
input	[15:0]	bus_51ae933d_;
input		bus_6a8dff02_;
input	[15:0]	bus_733d2b23_;
output	[15:0]	bus_70ada90a_;
wire		or_645c218d_u0;
reg	[15:0]	stateVar_rowRepeated_u3=16'h1;
wire	[15:0]	mux_4415bbea_u0;
wire	[15:0]	endianswapper_6acb6654_out;
wire	[15:0]	endianswapper_34cf1120_out;
assign or_645c218d_u0=bus_0469fc4f_|bus_6a8dff02_;
assign bus_70ada90a_=endianswapper_34cf1120_out;
always @(posedge bus_1d013d35_ or posedge bus_1beb5227_)
begin
if (bus_1beb5227_)
stateVar_rowRepeated_u3<=16'h1;
else if (or_645c218d_u0)
stateVar_rowRepeated_u3<=endianswapper_6acb6654_out;
end
assign mux_4415bbea_u0=(bus_0469fc4f_)?bus_51ae933d_:16'h1;
resized_LH1_xy_endianswapper_6acb6654_ resized_LH1_xy_endianswapper_6acb6654__1(.endianswapper_6acb6654_in(mux_4415bbea_u0), 
  .endianswapper_6acb6654_out(endianswapper_6acb6654_out));
resized_LH1_xy_endianswapper_34cf1120_ resized_LH1_xy_endianswapper_34cf1120__1(.endianswapper_34cf1120_in(stateVar_rowRepeated_u3), 
  .endianswapper_34cf1120_out(endianswapper_34cf1120_out));
endmodule



module resized_LH1_xy_structuralmemory_6d20861d_(CLK_u18, bus_28d40cb2_, bus_53538a8e_, bus_670f04d2_, bus_5f174387_, bus_3aeafa89_, bus_10b1614e_, bus_2d676b21_, bus_6bc2d2f4_);
input		CLK_u18;
input		bus_28d40cb2_;
input	[31:0]	bus_53538a8e_;
input	[2:0]	bus_670f04d2_;
input		bus_5f174387_;
input		bus_3aeafa89_;
input	[15:0]	bus_10b1614e_;
output	[15:0]	bus_2d676b21_;
output		bus_6bc2d2f4_;
wire		or_637c089e_u0;
reg		logicalMem_1e388226_we_delay0_u0=1'h0;
wire		or_20e47807_u0;
wire	[15:0]	bus_20a7b311_;
wire		and_4c630518_u0;
wire		not_215257c9_u0;
assign or_637c089e_u0=and_4c630518_u0|logicalMem_1e388226_we_delay0_u0;
always @(posedge CLK_u18 or posedge bus_28d40cb2_)
begin
if (bus_28d40cb2_)
logicalMem_1e388226_we_delay0_u0<=1'h0;
else logicalMem_1e388226_we_delay0_u0<=bus_3aeafa89_;
end
assign or_20e47807_u0=bus_5f174387_|bus_3aeafa89_;
assign bus_2d676b21_=bus_20a7b311_;
assign bus_6bc2d2f4_=or_637c089e_u0;
resized_LH1_xy_forge_memory_512x16_33 resized_LH1_xy_forge_memory_512x16_33_instance1(.CLK(CLK_u18), 
  .EN(or_20e47807_u0), .WE(bus_3aeafa89_), .ADDR(bus_53538a8e_), .DIN(bus_10b1614e_), 
  .DOUT(bus_20a7b311_), .DONE());
assign and_4c630518_u0=bus_5f174387_&not_215257c9_u0;
assign not_215257c9_u0=~bus_3aeafa89_;
endmodule



module resized_LH1_xy_consumeRow(CLK, RESET, GO, port_6e9d7dff_, port_2b507d31_, port_33a398fc_, port_58d4b229_, RESULT, RESULT_u1881, RESULT_u1882, RESULT_u1883, RESULT_u1884, RESULT_u1885, RESULT_u1886, RESULT_u1887, RESULT_u1888, RESULT_u1889, RESULT_u1890, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_6e9d7dff_;
input		port_2b507d31_;
input		port_33a398fc_;
input	[15:0]	port_58d4b229_;
output		RESULT;
output	[15:0]	RESULT_u1881;
output		RESULT_u1882;
output	[31:0]	RESULT_u1883;
output	[15:0]	RESULT_u1884;
output	[2:0]	RESULT_u1885;
output		RESULT_u1886;
output	[31:0]	RESULT_u1887;
output	[15:0]	RESULT_u1888;
output	[2:0]	RESULT_u1889;
output		RESULT_u1890;
output		DONE;
wire		simplePinWrite;
wire		and_u3173_u0;
wire		lessThanEqualTo;
wire signed	[16:0]	lessThanEqualTo_b_signed;
wire signed	[16:0]	lessThanEqualTo_a_signed;
wire		and_u3174_u0;
wire		not_u534_u0;
wire		and_u3175_u0;
reg		and_delayed_u214=1'h0;
wire	[31:0]	add;
wire	[31:0]	add_u375;
wire		or_u914_u0;
wire		and_u3176_u0;
reg		reg_2004ad98_u0=1'h0;
wire	[15:0]	add_u376;
reg	[15:0]	syncEnable_u559=16'h0;
wire		and_u3177_u0;
wire		or_u915_u0;
wire	[15:0]	mux_u335;
reg	[15:0]	latch_30329540_reg=16'h0;
wire	[15:0]	latch_30329540_out;
wire	[15:0]	add_u377;
wire		and_u3178_u0;
wire	[15:0]	subtract;
wire	[31:0]	add_u378;
wire		or_u916_u0;
wire		and_u3179_u0;
reg		reg_36fd5aa2_u0=1'h0;
wire	[15:0]	add_u379;
reg	[15:0]	syncEnable_u560_u0=16'h0;
wire signed	[16:0]	lessThanEqualTo_u3_b_signed;
wire		lessThanEqualTo_u3;
wire signed	[16:0]	lessThanEqualTo_u3_a_signed;
wire		not_u535_u0;
wire		and_u3180_u0;
wire		and_u3181_u0;
reg		reg_024cf124_u0=1'h0;
wire		and_u3182_u0;
reg	[15:0]	latch_47d885d0_reg=16'h0;
wire	[15:0]	latch_47d885d0_out;
wire		or_u917_u0;
wire	[15:0]	mux_u336_u0;
reg	[15:0]	syncEnable_u561_u0=16'h0;
reg		reg_1d7aa656_u0=1'h0;
assign simplePinWrite=GO&{1{GO}};
assign and_u3173_u0=and_u3174_u0&or_u915_u0;
assign lessThanEqualTo_a_signed={mux_u335[15], mux_u335};
assign lessThanEqualTo_b_signed=17'h1;
assign lessThanEqualTo=lessThanEqualTo_a_signed<=lessThanEqualTo_b_signed;
assign and_u3174_u0=or_u915_u0&lessThanEqualTo;
assign not_u534_u0=~lessThanEqualTo;
assign and_u3175_u0=or_u915_u0&not_u534_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u214<=1'h0;
else and_delayed_u214<=and_u3173_u0;
end
assign add={15'b0, port_6e9d7dff_, 1'b0}+{mux_u335[15], mux_u335[15], mux_u335[15], mux_u335[15], mux_u335[15], mux_u335[15], mux_u335[15], mux_u335[15], mux_u335[15], mux_u335[15], mux_u335[15], mux_u335[15], mux_u335[15], mux_u335[15], mux_u335[15], mux_u335[15], mux_u335};
assign add_u375={add[18], add[18], add[18], add[18], add[18], add[18], add[18], add[18], add[18], add[18], add[18], add[18], add[18], add[18:0]}+32'h0;
assign or_u914_u0=and_u3176_u0|RESET;
assign and_u3176_u0=reg_2004ad98_u0&port_2b507d31_;
always @(posedge CLK or posedge and_u3173_u0 or posedge or_u914_u0)
begin
if (or_u914_u0)
reg_2004ad98_u0<=1'h0;
else if (and_u3173_u0)
reg_2004ad98_u0<=1'h1;
else reg_2004ad98_u0<=reg_2004ad98_u0;
end
assign add_u376=mux_u335+16'h1;
always @(posedge CLK)
begin
if (and_u3173_u0)
syncEnable_u559<=add_u376;
end
assign and_u3177_u0=and_u3175_u0&or_u915_u0;
assign or_u915_u0=and_delayed_u214|GO;
assign mux_u335=(and_delayed_u214)?syncEnable_u559:16'h0;
always @(posedge CLK)
begin
if (GO)
latch_30329540_reg<=port_58d4b229_;
end
assign latch_30329540_out=(GO)?port_58d4b229_:latch_30329540_reg;
assign add_u377=port_6e9d7dff_+16'h1;
assign and_u3178_u0=and_u3181_u0&or_u917_u0;
assign subtract=mux_u336_u0-16'h1;
assign add_u378={subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract}+32'h0;
assign or_u916_u0=and_u3179_u0|RESET;
assign and_u3179_u0=reg_36fd5aa2_u0&port_33a398fc_;
always @(posedge CLK or posedge and_u3182_u0 or posedge or_u916_u0)
begin
if (or_u916_u0)
reg_36fd5aa2_u0<=1'h0;
else if (and_u3182_u0)
reg_36fd5aa2_u0<=1'h1;
else reg_36fd5aa2_u0<=reg_36fd5aa2_u0;
end
assign add_u379=mux_u336_u0+16'h1;
always @(posedge CLK)
begin
if (and_u3182_u0)
syncEnable_u560_u0<=add_u379;
end
assign lessThanEqualTo_u3_a_signed={mux_u336_u0[15], mux_u336_u0};
assign lessThanEqualTo_u3_b_signed=17'h2;
assign lessThanEqualTo_u3=lessThanEqualTo_u3_a_signed<=lessThanEqualTo_u3_b_signed;
assign not_u535_u0=~lessThanEqualTo_u3;
assign and_u3180_u0=or_u917_u0&lessThanEqualTo_u3;
assign and_u3181_u0=or_u917_u0&not_u535_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_024cf124_u0<=1'h0;
else reg_024cf124_u0<=and_u3182_u0;
end
assign and_u3182_u0=and_u3180_u0&or_u917_u0;
always @(posedge CLK)
begin
if (GO)
latch_47d885d0_reg<=port_58d4b229_;
end
assign latch_47d885d0_out=(GO)?port_58d4b229_:latch_47d885d0_reg;
assign or_u917_u0=reg_024cf124_u0|GO;
assign mux_u336_u0=(reg_024cf124_u0)?syncEnable_u560_u0:16'h1;
always @(posedge CLK)
begin
if (GO)
syncEnable_u561_u0<=add_u377;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1d7aa656_u0<=1'h0;
else reg_1d7aa656_u0<=and_u3177_u0;
end
assign RESULT=and_u3177_u0;
assign RESULT_u1881=syncEnable_u561_u0;
assign RESULT_u1882=and_u3173_u0;
assign RESULT_u1883=add_u375;
assign RESULT_u1884=latch_30329540_out;
assign RESULT_u1885=3'h1;
assign RESULT_u1886=and_u3182_u0;
assign RESULT_u1887=add_u378;
assign RESULT_u1888=latch_47d885d0_out;
assign RESULT_u1889=3'h1;
assign RESULT_u1890=simplePinWrite;
assign DONE=reg_1d7aa656_u0;
endmodule


