// __  ___ __ ___  _ __   ___  ___ 
// \ \/ / '__/ _ \| '_ \ / _ \/ __|
//  >  <| | | (_) | | | | (_) \__ \
// /_/\_\_|  \___/|_| |_|\___/|___/
// 
// Xronos synthesizer version
// Run date: Thu 2 Nov 2017 13:58:36 +0000
// 

module LL2_iunzip(In1_ACK, Out1_COUNT, Out2_DATA, CLK, RESET, Out1_SEND, In1_SEND, Out1_RDY, In1_COUNT, Out2_ACK, Out2_COUNT, In1_DATA, Out1_ACK, Out2_SEND, Out2_RDY, Out1_DATA);
wire		firstNPixels_done;
output		In1_ACK;
output	[15:0]	Out1_COUNT;
wire		streamEndFun1_done;
output	[15:0]	Out2_DATA;
wire		firstNPixels_go;
wire		streamEndFun2_go;
wire		streamEndFun2_done;
input		CLK;
input		RESET;
output		Out1_SEND;
wire		streamFun1_done;
wire		streamFun2_done;
input		In1_SEND;
input		Out1_RDY;
input	[15:0]	In1_COUNT;
input		Out2_ACK;
output	[15:0]	Out2_COUNT;
input	[15:0]	In1_DATA;
wire		streamFun1_go;
wire		streamFun2_go;
input		Out1_ACK;
output		Out2_SEND;
wire		streamEndFun1_go;
input		Out2_RDY;
output	[15:0]	Out1_DATA;
wire		bus_00559d40_;
wire		or_32361cb4_u0;
wire		bus_1f37da69_;
wire		bus_2d01cb3b_;
wire	[31:0]	bus_64537cfa_;
wire	[2:0]	bus_08021ab3_;
wire	[15:0]	bus_563cdce1_;
wire		bus_1dcb6638_;
wire		bus_23a30334_;
wire	[15:0]	bus_5e9e7e89_;
wire	[15:0]	bus_6317e79e_;
wire		bus_071890d3_;
wire	[15:0]	bus_3459005e_;
wire		bus_401a25a2_;
wire		bus_07cbf505_;
wire		or_6cb6ea2f_u0;
wire		streamEndFun1_u30;
wire		streamEndFun1_u26;
wire	[15:0]	streamEndFun1_u34;
wire	[15:0]	streamEndFun1_u33;
wire	[15:0]	streamEndFun1_u38;
wire	[2:0]	streamEndFun1_u29;
wire	[15:0]	streamEndFun1_u37;
wire	[31:0]	streamEndFun1_u31;
wire		streamEndFun1_u36;
wire		streamEndFun1_u27;
wire		streamEndFun1;
wire	[31:0]	streamEndFun1_u28;
wire		LL2_iunzip_streamEndFun1_instance_DONE;
wire	[2:0]	streamEndFun1_u32;
wire		streamEndFun1_u35;
wire	[31:0]	bus_32c38fb2_;
wire	[15:0]	or_718ad8aa_u0;
wire	[31:0]	bus_0e817a69_;
wire		bus_0c3d5734_;
wire	[1:0]	bus_3c983ce7_;
wire	[31:0]	bus_13fc03a5_;
wire		bus_09dd7fc4_;
wire		streamEndFun2_u30;
wire		streamEndFun2_u26;
wire	[31:0]	streamEndFun2_u31;
wire	[2:0]	streamEndFun2_u32;
wire	[15:0]	streamEndFun2_u33;
wire	[15:0]	streamEndFun2_u38;
wire	[15:0]	streamEndFun2_u37;
wire		streamEndFun2_u27;
wire	[15:0]	streamEndFun2_u34;
wire		LL2_iunzip_streamEndFun2_instance_DONE;
wire	[31:0]	streamEndFun2_u28;
wire		streamEndFun2;
wire		streamEndFun2_u36;
wire		streamEndFun2_u35;
wire	[2:0]	streamEndFun2_u29;
wire	[1:0]	bus_3078af4b_;
wire	[2:0]	streamFun2_u43;
wire	[2:0]	streamFun2_u40;
wire	[2:0]	streamFun2_u46;
wire		streamFun2_u41;
wire		streamFun2_u35;
wire		streamFun2;
wire		streamFun2_u48;
wire		streamFun2_u44;
wire		streamFun2_u37;
wire		streamFun2_u49;
wire	[31:0]	streamFun2_u36;
wire	[15:0]	streamFun2_u50;
wire	[31:0]	streamFun2_u45;
wire	[31:0]	streamFun2_u38;
wire	[15:0]	streamFun2_u39;
wire		LL2_iunzip_streamFun2_instance_DONE;
wire	[15:0]	streamFun2_u47;
wire	[31:0]	streamFun2_u42;
wire		streamFun2_u34;
wire	[31:0]	bus_1d7ad841_;
wire		bus_1d3acc5f_;
wire	[15:0]	bus_6715655d_;
wire		bus_36f7a4bd_;
wire	[2:0]	bus_7046b040_;
wire	[15:0]	bus_005f3f40_;
wire		bus_6d1b31d9_;
wire	[15:0]	or_235a4690_u0;
wire	[15:0]	or_14287ce5_u0;
wire		bus_0c01b8a2_;
wire	[15:0]	bus_29133072_;
wire		bus_52940f8a_;
wire	[15:0]	bus_066c060a_;
wire		bus_7c6d4762_;
wire		bus_01050093_;
wire		bus_7db96305_;
wire	[2:0]	bus_79309e44_;
wire	[15:0]	bus_5a3ab128_;
wire		bus_539df49f_;
wire	[15:0]	bus_7e0b6b8d_;
wire	[15:0]	bus_5263a0f6_;
wire	[15:0]	bus_7045541b_;
wire	[31:0]	bus_2873baa2_;
wire		bus_72817d63_;
wire		bus_0e4c9451_;
wire		bus_44703396_;
wire	[15:0]	bus_7ca96f1c_;
wire		bus_7cd847a6_;
wire		scheduler_u145;
wire	[1:0]	scheduler_u138;
wire		LL2_iunzip_scheduler_instance_DONE;
wire		scheduler_u151;
wire	[31:0]	scheduler_u140;
wire	[31:0]	scheduler_u146;
wire		scheduler;
wire		scheduler_u139;
wire		scheduler_u144;
wire		scheduler_u149;
wire		scheduler_u150;
wire		scheduler_u153;
wire		scheduler_u152;
wire		scheduler_u143;
wire		scheduler_u137;
wire	[31:0]	scheduler_u142;
wire	[15:0]	scheduler_u147;
wire	[1:0]	scheduler_u136;
wire		scheduler_u141;
wire		scheduler_u154;
wire	[2:0]	scheduler_u148;
wire		bus_6ac01b98_;
wire	[15:0]	or_529e2dc5_u0;
wire		bus_60f9b471_;
wire		or_06358b68_u0;
wire	[15:0]	bus_5ab9ae07_;
wire	[2:0]	bus_7e94d1e2_;
wire		bus_1c0ab1f7_;
wire		bus_4174f34a_;
wire		bus_1b8550b0_;
wire	[15:0]	bus_0a857fee_;
wire	[15:0]	bus_51d68f43_;
wire		bus_0e2119bf_;
wire	[15:0]	bus_22cdc0fd_;
wire		bus_33af47da_;
wire	[31:0]	bus_3266894e_;
wire	[15:0]	bus_098f7792_;
wire		bus_49128048_;
wire		bus_38e1176c_;
wire		streamFun1_u48;
wire	[2:0]	streamFun1_u43;
wire	[31:0]	streamFun1_u45;
wire		streamFun1_u35;
wire	[2:0]	streamFun1_u39;
wire		streamFun1_u44;
wire	[15:0]	streamFun1_u50;
wire		streamFun1;
wire		streamFun1_u34;
wire	[31:0]	streamFun1_u36;
wire		streamFun1_u49;
wire	[31:0]	streamFun1_u38;
wire	[15:0]	streamFun1_u42;
wire	[15:0]	streamFun1_u47;
wire		streamFun1_u40;
wire		LL2_iunzip_streamFun1_instance_DONE;
wire		streamFun1_u37;
wire	[31:0]	streamFun1_u41;
wire	[2:0]	streamFun1_u46;
wire		firstNPixels_u23;
wire	[31:0]	firstNPixels_u31;
wire		firstNPixels;
wire	[2:0]	firstNPixels_u25;
wire		LL2_iunzip_firstNPixels_instance_DONE;
wire		firstNPixels_u26;
wire	[31:0]	firstNPixels_u22;
wire	[2:0]	firstNPixels_u29;
wire	[2:0]	firstNPixels_u32;
wire	[31:0]	firstNPixels_u27;
wire		firstNPixels_u30;
wire	[31:0]	firstNPixels_u24;
wire	[15:0]	firstNPixels_u28;
wire		bus_137455cf_;
assign firstNPixels_done=bus_09dd7fc4_;
assign In1_ACK=or_6cb6ea2f_u0;
assign Out1_COUNT=or_235a4690_u0;
assign streamEndFun1_done=bus_0c3d5734_;
assign Out2_DATA=or_718ad8aa_u0;
assign firstNPixels_go=scheduler_u153;
assign streamEndFun2_go=scheduler_u149;
assign streamEndFun2_done=bus_00559d40_;
assign Out1_SEND=or_32361cb4_u0;
assign streamFun1_done=bus_7cd847a6_;
assign streamFun2_done=bus_60f9b471_;
assign Out2_COUNT=or_529e2dc5_u0;
assign streamFun1_go=scheduler_u150;
assign streamFun2_go=scheduler_u151;
assign Out2_SEND=or_06358b68_u0;
assign streamEndFun1_go=scheduler_u154;
assign Out1_DATA=or_14287ce5_u0;
assign bus_00559d40_=LL2_iunzip_streamEndFun2_instance_DONE&{1{LL2_iunzip_streamEndFun2_instance_DONE}};
assign or_32361cb4_u0=streamFun1_u48|streamEndFun1_u35|streamEndFun2_u35;
LL2_iunzip_simplememoryreferee_2945e249_ LL2_iunzip_simplememoryreferee_2945e249__1(.bus_2951946e_(CLK), 
  .bus_416e1391_(bus_38e1176c_), .bus_2a47c7a6_(bus_0c01b8a2_), .bus_7242c66a_(bus_066c060a_), 
  .bus_4e73801e_(firstNPixels_u30), .bus_0e6b979a_(32'h0), .bus_15f2220c_(3'h1), 
  .bus_71d990b7_(scheduler_u145), .bus_0fb935b7_(scheduler_u147), .bus_3e195330_(scheduler_u146), 
  .bus_61a7ee67_(3'h1), .bus_5e9e7e89_(bus_5e9e7e89_), .bus_64537cfa_(bus_64537cfa_), 
  .bus_2d01cb3b_(bus_2d01cb3b_), .bus_1f37da69_(bus_1f37da69_), .bus_08021ab3_(bus_08021ab3_), 
  .bus_563cdce1_(bus_563cdce1_), .bus_1dcb6638_(bus_1dcb6638_), .bus_23a30334_(bus_23a30334_));
LL2_iunzip_structuralmemory_0dd5b544_ LL2_iunzip_structuralmemory_0dd5b544__1(.CLK_u6(CLK), 
  .bus_6e2d8210_(bus_38e1176c_), .bus_0cec7947_(bus_3266894e_), .bus_0faf4bd2_(3'h1), 
  .bus_675a5739_(bus_1b8550b0_), .bus_7124b784_(bus_2873baa2_), .bus_12baf768_(3'h1), 
  .bus_1b5dd815_(bus_7c6d4762_), .bus_45524d51_(bus_7db96305_), .bus_25748481_(bus_7ca96f1c_), 
  .bus_6317e79e_(bus_6317e79e_), .bus_071890d3_(bus_071890d3_), .bus_3459005e_(bus_3459005e_), 
  .bus_401a25a2_(bus_401a25a2_));
LL2_iunzip_Kicker_30 LL2_iunzip_Kicker_30_1(.CLK(CLK), .RESET(bus_38e1176c_), .bus_07cbf505_(bus_07cbf505_));
assign or_6cb6ea2f_u0=streamFun1_u49|streamFun2_u49|scheduler_u152;
LL2_iunzip_streamEndFun1 LL2_iunzip_streamEndFun1_instance(.CLK(CLK), .RESET(bus_38e1176c_), 
  .GO(streamEndFun1_go), .port_27264123_(bus_137455cf_), .port_20d55f53_(bus_539df49f_), 
  .port_0a0c52a4_(bus_7045541b_), .port_2c516464_(bus_33af47da_), .port_5613faef_(bus_22cdc0fd_), 
  .DONE(LL2_iunzip_streamEndFun1_instance_DONE), .RESULT(streamEndFun1), .RESULT_u950(streamEndFun1_u26), 
  .RESULT_u954(streamEndFun1_u27), .RESULT_u955(streamEndFun1_u28), .RESULT_u956(streamEndFun1_u29), 
  .RESULT_u951(streamEndFun1_u30), .RESULT_u952(streamEndFun1_u31), .RESULT_u953(streamEndFun1_u32), 
  .RESULT_u957(streamEndFun1_u33), .RESULT_u958(streamEndFun1_u34), .RESULT_u959(streamEndFun1_u35), 
  .RESULT_u960(streamEndFun1_u36), .RESULT_u961(streamEndFun1_u37), .RESULT_u962(streamEndFun1_u38));
LL2_iunzip_stateVar_In1TokenIndex LL2_iunzip_stateVar_In1TokenIndex_1(.bus_221c1ac8_(CLK), 
  .bus_4e95ce1d_(bus_38e1176c_), .bus_119618fb_(scheduler_u139), .bus_339b4303_(scheduler_u140), 
  .bus_32c38fb2_(bus_32c38fb2_));
assign or_718ad8aa_u0=streamFun2_u50|streamEndFun1_u38|streamEndFun2_u38;
LL2_iunzip_stateVar_In1MaxTokenIndex LL2_iunzip_stateVar_In1MaxTokenIndex_1(.bus_54c26aa4_(CLK), 
  .bus_19793f6e_(bus_38e1176c_), .bus_299324f7_(scheduler_u141), .bus_3e112cd2_({scheduler_u142[31:2], 1'b0, scheduler_u142[0]}), 
  .bus_0e817a69_(bus_0e817a69_));
assign bus_0c3d5734_=LL2_iunzip_streamEndFun1_instance_DONE&{1{LL2_iunzip_streamEndFun1_instance_DONE}};
LL2_iunzip_stateVar_fsmState_LL2_iunzip LL2_iunzip_stateVar_fsmState_LL2_iunzip_1(.bus_2d067e63_(CLK), 
  .bus_38ab1e34_(bus_38e1176c_), .bus_3d48ec63_(scheduler_u137), .bus_43199831_(scheduler_u138), 
  .bus_3c983ce7_(bus_3c983ce7_));
LL2_iunzip_stateVar_consumed LL2_iunzip_stateVar_consumed_1(.bus_416e1293_(CLK), 
  .bus_12087713_(bus_38e1176c_), .bus_191cf97c_(firstNPixels), .bus_79b6c0b0_(firstNPixels_u22), 
  .bus_3df41d15_(streamFun1_u35), .bus_6619539b_(streamFun1_u36), .bus_5630e916_(streamFun2_u35), 
  .bus_7ed235d5_(streamFun2_u36), .bus_13fc03a5_(bus_13fc03a5_));
assign bus_09dd7fc4_=LL2_iunzip_firstNPixels_instance_DONE&{1{LL2_iunzip_firstNPixels_instance_DONE}};
LL2_iunzip_streamEndFun2 LL2_iunzip_streamEndFun2_instance(.CLK(CLK), .RESET(bus_38e1176c_), 
  .GO(streamEndFun2_go), .port_2a8e19bd_(bus_137455cf_), .port_377c7b5e_(bus_0e2119bf_), 
  .port_3606eb83_(bus_51d68f43_), .port_1d8d2ce2_(bus_0e4c9451_), .port_2bdba753_(bus_5263a0f6_), 
  .DONE(LL2_iunzip_streamEndFun2_instance_DONE), .RESULT(streamEndFun2), .RESULT_u963(streamEndFun2_u26), 
  .RESULT_u964(streamEndFun2_u27), .RESULT_u965(streamEndFun2_u28), .RESULT_u966(streamEndFun2_u29), 
  .RESULT_u967(streamEndFun2_u30), .RESULT_u968(streamEndFun2_u31), .RESULT_u969(streamEndFun2_u32), 
  .RESULT_u970(streamEndFun2_u33), .RESULT_u971(streamEndFun2_u34), .RESULT_u972(streamEndFun2_u35), 
  .RESULT_u973(streamEndFun2_u36), .RESULT_u974(streamEndFun2_u37), .RESULT_u975(streamEndFun2_u38));
LL2_iunzip_stateVar_fsmOldState_LL2_iunzip LL2_iunzip_stateVar_fsmOldState_LL2_iunzip_1(.bus_3b581e33_(CLK), 
  .bus_52d5710c_(bus_38e1176c_), .bus_4ec3c878_(scheduler), .bus_4cb5a4aa_(scheduler_u136), 
  .bus_3078af4b_(bus_3078af4b_));
LL2_iunzip_streamFun2 LL2_iunzip_streamFun2_instance(.CLK(CLK), .RESET(bus_38e1176c_), 
  .GO(streamFun2_go), .port_5fca059d_(bus_137455cf_), .port_581d88d1_(bus_13fc03a5_), 
  .port_4ccd3ea3_(bus_44703396_), .port_79fe3347_(bus_1c0ab1f7_), .port_3b68465d_(bus_098f7792_), 
  .port_7396b25e_(bus_44703396_), .port_33e93e76_(bus_7e0b6b8d_), .port_2d7037ba_(In1_DATA), 
  .DONE(LL2_iunzip_streamFun2_instance_DONE), .RESULT(streamFun2), .RESULT_u976(streamFun2_u34), 
  .RESULT_u977(streamFun2_u35), .RESULT_u978(streamFun2_u36), .RESULT_u985(streamFun2_u37), 
  .RESULT_u986(streamFun2_u38), .RESULT_u987(streamFun2_u39), .RESULT_u988(streamFun2_u40), 
  .RESULT_u979(streamFun2_u41), .RESULT_u980(streamFun2_u42), .RESULT_u981(streamFun2_u43), 
  .RESULT_u982(streamFun2_u44), .RESULT_u983(streamFun2_u45), .RESULT_u984(streamFun2_u46), 
  .RESULT_u989(streamFun2_u47), .RESULT_u990(streamFun2_u48), .RESULT_u991(streamFun2_u49), 
  .RESULT_u992(streamFun2_u50));
LL2_iunzip_simplememoryreferee_15caad00_ LL2_iunzip_simplememoryreferee_15caad00__1(.bus_16cdabb7_(CLK), 
  .bus_0de57dc4_(bus_38e1176c_), .bus_7b32a18c_(bus_52940f8a_), .bus_247edfb6_(bus_29133072_), 
  .bus_229405ff_(firstNPixels_u23), .bus_5a473665_(32'h1), .bus_36b4444a_(3'h1), 
  .bus_005f3f40_(bus_005f3f40_), .bus_1d7ad841_(bus_1d7ad841_), .bus_36f7a4bd_(bus_36f7a4bd_), 
  .bus_6d1b31d9_(bus_6d1b31d9_), .bus_7046b040_(bus_7046b040_), .bus_6715655d_(bus_6715655d_), 
  .bus_1d3acc5f_(bus_1d3acc5f_));
assign or_235a4690_u0=streamFun1_u50|streamEndFun1_u37|streamEndFun2_u37;
assign or_14287ce5_u0=streamFun1_u47|streamEndFun1_u34|streamEndFun2_u34;
LL2_iunzip_structuralmemory_0e000751_ LL2_iunzip_structuralmemory_0e000751__1(.CLK_u7(CLK), 
  .bus_457d065b_(bus_38e1176c_), .bus_417f17f6_(32'h1), .bus_7399bd45_(3'h1), .bus_6a7bbc81_(bus_6d1b31d9_), 
  .bus_3cbe9f79_(bus_64537cfa_), .bus_04ea2051_(3'h1), .bus_4640c3a2_(bus_1f37da69_), 
  .bus_73e3f3e7_(bus_2d01cb3b_), .bus_4ce023f4_(bus_5e9e7e89_), .bus_29133072_(bus_29133072_), 
  .bus_52940f8a_(bus_52940f8a_), .bus_066c060a_(bus_066c060a_), .bus_0c01b8a2_(bus_0c01b8a2_));
LL2_iunzip_simplememoryreferee_06e2d637_ LL2_iunzip_simplememoryreferee_06e2d637__1(.bus_54a19bc9_(CLK), 
  .bus_4453c8b0_(bus_38e1176c_), .bus_567d4ed5_(bus_401a25a2_), .bus_59677524_(bus_3459005e_), 
  .bus_209bc1d3_(firstNPixels_u26), .bus_2383042c_(firstNPixels_u28), .bus_355229bb_({31'b0, firstNPixels_u27[0]}), 
  .bus_765ef4b2_(3'h1), .bus_23a9aa5b_(streamFun1_u37), .bus_0d9a64c8_(streamFun1_u40), 
  .bus_17a89a93_(streamFun1_u42), .bus_5555630d_(streamFun1_u41), .bus_3552a76c_(3'h1), 
  .bus_57a3f872_(streamFun2_u44), .bus_5ee3d6e0_(streamFun2_u37), .bus_6483aa66_(streamFun2_u39), 
  .bus_6cf5cfbb_(streamFun2_u38), .bus_62f7ce09_(3'h1), .bus_35ec3db3_(streamEndFun1_u27), 
  .bus_27b331c3_(streamEndFun1_u28), .bus_14e11e79_(3'h1), .bus_6ee688b9_(streamEndFun2_u30), 
  .bus_2284bbc7_(streamEndFun2_u31), .bus_1c9a0cac_(3'h1), .bus_7ca96f1c_(bus_7ca96f1c_), 
  .bus_2873baa2_(bus_2873baa2_), .bus_7db96305_(bus_7db96305_), .bus_7c6d4762_(bus_7c6d4762_), 
  .bus_79309e44_(bus_79309e44_), .bus_72817d63_(bus_72817d63_), .bus_5a3ab128_(bus_5a3ab128_), 
  .bus_01050093_(bus_01050093_), .bus_7e0b6b8d_(bus_7e0b6b8d_), .bus_44703396_(bus_44703396_), 
  .bus_7045541b_(bus_7045541b_), .bus_539df49f_(bus_539df49f_), .bus_5263a0f6_(bus_5263a0f6_), 
  .bus_0e4c9451_(bus_0e4c9451_));
assign bus_7cd847a6_=LL2_iunzip_streamFun1_instance_DONE&{1{LL2_iunzip_streamFun1_instance_DONE}};
LL2_iunzip_scheduler LL2_iunzip_scheduler_instance(.CLK(CLK), .RESET(bus_38e1176c_), 
  .GO(bus_07cbf505_), .port_44cbc7ff_(bus_3078af4b_), .port_57df124f_(bus_3c983ce7_), 
  .port_2710208c_(bus_32c38fb2_), .port_0dedb00e_(bus_0e817a69_), .port_0cb02262_(bus_13fc03a5_), 
  .port_51623660_(bus_23a30334_), .port_5f577b2f_(streamFun2_done), .port_2d918d8b_(In1_SEND), 
  .port_3777dab3_(Out2_RDY), .port_6a679525_(streamEndFun2_done), .port_5a872d3c_(In1_DATA), 
  .port_1a1203bd_(firstNPixels_done), .port_4cbbb047_(Out1_RDY), .port_59e64907_(streamEndFun1_done), 
  .port_5351796d_(streamFun1_done), .DONE(LL2_iunzip_scheduler_instance_DONE), 
  .RESULT(scheduler), .RESULT_u993(scheduler_u136), .RESULT_u994(scheduler_u137), 
  .RESULT_u995(scheduler_u138), .RESULT_u996(scheduler_u139), .RESULT_u997(scheduler_u140), 
  .RESULT_u998(scheduler_u141), .RESULT_u999(scheduler_u142), .RESULT_u1000(scheduler_u143), 
  .RESULT_u1001(scheduler_u144), .RESULT_u1002(scheduler_u145), .RESULT_u1003(scheduler_u146), 
  .RESULT_u1004(scheduler_u147), .RESULT_u1005(scheduler_u148), .RESULT_u1006(scheduler_u149), 
  .RESULT_u1007(scheduler_u150), .RESULT_u1008(scheduler_u151), .RESULT_u1009(scheduler_u152), 
  .RESULT_u1010(scheduler_u153), .RESULT_u1011(scheduler_u154));
LL2_iunzip_stateVar_In1PortEnable LL2_iunzip_stateVar_In1PortEnable_1(.bus_4b677821_(CLK), 
  .bus_30c4b424_(bus_38e1176c_), .bus_2657c6ba_(scheduler_u143), .bus_4371ff51_(scheduler_u144), 
  .bus_6ac01b98_(bus_6ac01b98_));
assign or_529e2dc5_u0=streamFun2_u47|streamEndFun1_u33|streamEndFun2_u33;
assign bus_60f9b471_=LL2_iunzip_streamFun2_instance_DONE&{1{LL2_iunzip_streamFun2_instance_DONE}};
assign or_06358b68_u0=streamFun2_u48|streamEndFun1_u36|streamEndFun2_u36;
LL2_iunzip_simplememoryreferee_27761197_ LL2_iunzip_simplememoryreferee_27761197__1(.bus_60b63314_(CLK), 
  .bus_0869b5ee_(bus_38e1176c_), .bus_764c86ba_(bus_071890d3_), .bus_43e4e98d_(bus_6317e79e_), 
  .bus_52c6af95_(streamFun1_u44), .bus_524a4e4b_(streamFun1_u45), .bus_43a489ea_(3'h1), 
  .bus_5442bd92_(streamFun2_u41), .bus_1328384d_(streamFun2_u42), .bus_73af1459_(3'h1), 
  .bus_6b014163_(streamEndFun1_u30), .bus_4135f178_(streamEndFun1_u31), .bus_6616c9bf_(3'h1), 
  .bus_188e8a1f_(streamEndFun2_u27), .bus_79e17b19_(streamEndFun2_u28), .bus_055751fe_(3'h1), 
  .bus_5ab9ae07_(bus_5ab9ae07_), .bus_3266894e_(bus_3266894e_), .bus_4174f34a_(bus_4174f34a_), 
  .bus_1b8550b0_(bus_1b8550b0_), .bus_7e94d1e2_(bus_7e94d1e2_), .bus_0a857fee_(bus_0a857fee_), 
  .bus_49128048_(bus_49128048_), .bus_098f7792_(bus_098f7792_), .bus_1c0ab1f7_(bus_1c0ab1f7_), 
  .bus_22cdc0fd_(bus_22cdc0fd_), .bus_33af47da_(bus_33af47da_), .bus_51d68f43_(bus_51d68f43_), 
  .bus_0e2119bf_(bus_0e2119bf_));
LL2_iunzip_globalreset_physical_4d3e90cc_ LL2_iunzip_globalreset_physical_4d3e90cc__1(.bus_7a7df9cf_(CLK), 
  .bus_50fc0f9a_(RESET), .bus_38e1176c_(bus_38e1176c_));
LL2_iunzip_streamFun1 LL2_iunzip_streamFun1_instance(.CLK(CLK), .RESET(bus_38e1176c_), 
  .GO(streamFun1_go), .port_02b645ca_(bus_137455cf_), .port_782b7e63_(bus_13fc03a5_), 
  .port_45c60a90_(bus_01050093_), .port_02d3b259_(bus_5a3ab128_), .port_73617117_(bus_01050093_), 
  .port_678d8025_(bus_49128048_), .port_6a7883c4_(bus_0a857fee_), .port_32d96ef1_(In1_DATA), 
  .DONE(LL2_iunzip_streamFun1_instance_DONE), .RESULT(streamFun1), .RESULT_u1012(streamFun1_u34), 
  .RESULT_u1013(streamFun1_u35), .RESULT_u1014(streamFun1_u36), .RESULT_u1018(streamFun1_u37), 
  .RESULT_u1019(streamFun1_u38), .RESULT_u1020(streamFun1_u39), .RESULT_u1021(streamFun1_u40), 
  .RESULT_u1022(streamFun1_u41), .RESULT_u1023(streamFun1_u42), .RESULT_u1024(streamFun1_u43), 
  .RESULT_u1015(streamFun1_u44), .RESULT_u1016(streamFun1_u45), .RESULT_u1017(streamFun1_u46), 
  .RESULT_u1025(streamFun1_u47), .RESULT_u1026(streamFun1_u48), .RESULT_u1027(streamFun1_u49), 
  .RESULT_u1028(streamFun1_u50));
LL2_iunzip_firstNPixels LL2_iunzip_firstNPixels_instance(.CLK(CLK), .RESET(bus_38e1176c_), 
  .GO(firstNPixels_go), .port_56c10d09_(bus_13fc03a5_), .port_4bf45ad9_(bus_1d3acc5f_), 
  .port_5d69d1a2_(bus_6715655d_), .port_4285ced0_(bus_72817d63_), .port_7e889a85_(bus_1dcb6638_), 
  .port_7d5897f1_(bus_563cdce1_), .DONE(LL2_iunzip_firstNPixels_instance_DONE), 
  .RESULT(firstNPixels), .RESULT_u1029(firstNPixels_u22), .RESULT_u1037(firstNPixels_u23), 
  .RESULT_u1038(firstNPixels_u24), .RESULT_u1039(firstNPixels_u25), .RESULT_u1030(firstNPixels_u26), 
  .RESULT_u1031(firstNPixels_u27), .RESULT_u1032(firstNPixels_u28), .RESULT_u1033(firstNPixels_u29), 
  .RESULT_u1034(firstNPixels_u30), .RESULT_u1035(firstNPixels_u31), .RESULT_u1036(firstNPixels_u32));
LL2_iunzip_stateVar_midPoint LL2_iunzip_stateVar_midPoint_1(.bus_68e44dca_(CLK), 
  .bus_1d3a1112_(bus_38e1176c_), .bus_0b5520fb_(streamFun1), .bus_0cea9df7_(1'h0), 
  .bus_37b6d949_(streamFun2), .bus_03a0d5c2_(1'h0), .bus_24329444_(streamEndFun1), 
  .bus_150341ad_(1'h0), .bus_7bdb1d62_(streamEndFun2), .bus_20c3ad1e_(1'h0), .bus_137455cf_(bus_137455cf_));
endmodule



module LL2_iunzip_simplememoryreferee_2945e249_(bus_2951946e_, bus_416e1391_, bus_2a47c7a6_, bus_7242c66a_, bus_4e73801e_, bus_0e6b979a_, bus_15f2220c_, bus_71d990b7_, bus_0fb935b7_, bus_3e195330_, bus_61a7ee67_, bus_5e9e7e89_, bus_64537cfa_, bus_2d01cb3b_, bus_1f37da69_, bus_08021ab3_, bus_563cdce1_, bus_1dcb6638_, bus_23a30334_);
input		bus_2951946e_;
input		bus_416e1391_;
input		bus_2a47c7a6_;
input	[15:0]	bus_7242c66a_;
input		bus_4e73801e_;
input	[31:0]	bus_0e6b979a_;
input	[2:0]	bus_15f2220c_;
input		bus_71d990b7_;
input	[15:0]	bus_0fb935b7_;
input	[31:0]	bus_3e195330_;
input	[2:0]	bus_61a7ee67_;
output	[15:0]	bus_5e9e7e89_;
output	[31:0]	bus_64537cfa_;
output		bus_2d01cb3b_;
output		bus_1f37da69_;
output	[2:0]	bus_08021ab3_;
output	[15:0]	bus_563cdce1_;
output		bus_1dcb6638_;
output		bus_23a30334_;
wire		or_244305e6_u0;
reg		done_qual_u64=1'h0;
wire		or_2e648e2d_u0;
wire	[15:0]	mux_5bb34d01_u0;
wire	[31:0]	mux_68d17742_u0;
wire		or_70c06e94_u0;
wire		and_6833d967_u0;
wire		not_7393cc44_u0;
wire		not_0b3493e8_u0;
reg		done_qual_u65_u0=1'h0;
wire		and_58d64e49_u0;
assign bus_5e9e7e89_=mux_5bb34d01_u0;
assign bus_64537cfa_=mux_68d17742_u0;
assign bus_2d01cb3b_=bus_71d990b7_;
assign bus_1f37da69_=or_244305e6_u0;
assign bus_08021ab3_=3'h1;
assign bus_563cdce1_=bus_7242c66a_;
assign bus_1dcb6638_=and_58d64e49_u0;
assign bus_23a30334_=and_6833d967_u0;
assign or_244305e6_u0=bus_4e73801e_|bus_71d990b7_;
always @(posedge bus_2951946e_)
begin
if (bus_416e1391_)
done_qual_u64<=1'h0;
else done_qual_u64<=bus_4e73801e_;
end
assign or_2e648e2d_u0=bus_71d990b7_|done_qual_u65_u0;
assign mux_5bb34d01_u0=({16{bus_71d990b7_}}&bus_0fb935b7_);
assign mux_68d17742_u0=(bus_4e73801e_)?32'h0:bus_3e195330_;
assign or_70c06e94_u0=bus_4e73801e_|done_qual_u64;
assign and_6833d967_u0=or_2e648e2d_u0&bus_2a47c7a6_;
assign not_7393cc44_u0=~bus_2a47c7a6_;
assign not_0b3493e8_u0=~bus_2a47c7a6_;
always @(posedge bus_2951946e_)
begin
if (bus_416e1391_)
done_qual_u65_u0<=1'h0;
else done_qual_u65_u0<=bus_71d990b7_;
end
assign and_58d64e49_u0=or_70c06e94_u0&bus_2a47c7a6_;
endmodule



module LL2_iunzip_forge_memory_3x16_14(CLK, ENA, WEA, DINA, ENB, ADDRA, ADDRB, DOUTA, DOUTB, DONEA, DONEB);
input		CLK;
input		ENA;
input		WEA;
input	[15:0]	DINA;
input		ENB;
input	[31:0]	ADDRA;
input	[31:0]	ADDRB;
output	[15:0]	DOUTA;
output	[15:0]	DOUTB;
output		DONEA;
output		DONEB;
wire		wea_0;
wire	[15:0]	pre_douta_0;
wire	[15:0]	pre_doutb_0;
reg		wea_done;
reg		rea_done;
reg	[15:0]	mux_outa;
reg	[15:0]	mux_outb;
assign wea_0=WEA;
always @(posedge CLK)
begin
wea_done<=WEA;
end
assign DONEA=rea_done|wea_done;
always @(posedge CLK)
begin
end
assign DONEB=ENB;
always @(pre_douta_0)
begin
mux_outa<=pre_douta_0;
end
assign DOUTA=mux_outa;
always @(pre_doutb_0)
begin
mux_outb<=pre_doutb_0;
end
assign DOUTB=mux_outb;
// Memory array element: COL: 0, ROW: 0
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_64(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[0]), .SPO(pre_douta_0[0]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[0]));
// Memory array element: COL: 0, ROW: 1
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_65(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[1]), .SPO(pre_douta_0[1]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[1]));
// Memory array element: COL: 0, ROW: 2
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_66(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[2]), .SPO(pre_douta_0[2]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[2]));
// Memory array element: COL: 0, ROW: 3
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_67(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[3]), .SPO(pre_douta_0[3]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[3]));
// Memory array element: COL: 0, ROW: 4
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_68(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[4]), .SPO(pre_douta_0[4]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[4]));
// Memory array element: COL: 0, ROW: 5
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_69(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[5]), .SPO(pre_douta_0[5]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[5]));
// Memory array element: COL: 0, ROW: 6
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_70(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[6]), .SPO(pre_douta_0[6]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[6]));
// Memory array element: COL: 0, ROW: 7
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_71(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[7]), .SPO(pre_douta_0[7]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[7]));
// Memory array element: COL: 0, ROW: 8
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_72(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[8]), .SPO(pre_douta_0[8]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[8]));
// Memory array element: COL: 0, ROW: 9
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_73(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[9]), .SPO(pre_douta_0[9]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[9]));
// Memory array element: COL: 0, ROW: 10
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_74(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[10]), .SPO(pre_douta_0[10]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[10]));
// Memory array element: COL: 0, ROW: 11
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_75(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[11]), .SPO(pre_douta_0[11]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[11]));
// Memory array element: COL: 0, ROW: 12
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_76(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[12]), .SPO(pre_douta_0[12]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[12]));
// Memory array element: COL: 0, ROW: 13
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_77(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[13]), .SPO(pre_douta_0[13]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[13]));
// Memory array element: COL: 0, ROW: 14
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_78(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[14]), .SPO(pre_douta_0[14]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[14]));
// Memory array element: COL: 0, ROW: 15
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_79(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[15]), .SPO(pre_douta_0[15]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[15]));
endmodule



module LL2_iunzip_structuralmemory_0dd5b544_(CLK_u6, bus_6e2d8210_, bus_0cec7947_, bus_0faf4bd2_, bus_675a5739_, bus_7124b784_, bus_12baf768_, bus_1b5dd815_, bus_45524d51_, bus_25748481_, bus_6317e79e_, bus_071890d3_, bus_3459005e_, bus_401a25a2_);
input		CLK_u6;
input		bus_6e2d8210_;
input	[31:0]	bus_0cec7947_;
input	[2:0]	bus_0faf4bd2_;
input		bus_675a5739_;
input	[31:0]	bus_7124b784_;
input	[2:0]	bus_12baf768_;
input		bus_1b5dd815_;
input		bus_45524d51_;
input	[15:0]	bus_25748481_;
output	[15:0]	bus_6317e79e_;
output		bus_071890d3_;
output	[15:0]	bus_3459005e_;
output		bus_401a25a2_;
wire		or_68602180_u0;
reg		logicalMem_74b878c1_we_delay0_u0=1'h0;
wire		and_0a1cb6b6_u0;
wire	[15:0]	bus_04c2aad9_;
wire	[15:0]	bus_0f2bbba2_;
wire		not_319421e2_u0;
wire		or_4c925a8c_u0;
assign or_68602180_u0=bus_1b5dd815_|bus_45524d51_;
always @(posedge CLK_u6 or posedge bus_6e2d8210_)
begin
if (bus_6e2d8210_)
logicalMem_74b878c1_we_delay0_u0<=1'h0;
else logicalMem_74b878c1_we_delay0_u0<=bus_45524d51_;
end
assign and_0a1cb6b6_u0=bus_1b5dd815_&not_319421e2_u0;
LL2_iunzip_forge_memory_3x16_14 LL2_iunzip_forge_memory_3x16_14_instance0(.CLK(CLK_u6), 
  .ENA(or_68602180_u0), .WEA(bus_45524d51_), .DINA(bus_25748481_), .ADDRA(bus_7124b784_), 
  .DOUTA(bus_04c2aad9_), .DONEA(), .ENB(bus_675a5739_), .ADDRB(bus_0cec7947_), .DOUTB(bus_0f2bbba2_), 
  .DONEB());
assign not_319421e2_u0=~bus_45524d51_;
assign bus_6317e79e_=bus_0f2bbba2_;
assign bus_071890d3_=bus_675a5739_;
assign bus_3459005e_=bus_04c2aad9_;
assign bus_401a25a2_=or_4c925a8c_u0;
assign or_4c925a8c_u0=and_0a1cb6b6_u0|logicalMem_74b878c1_we_delay0_u0;
endmodule



module LL2_iunzip_Kicker_30(CLK, RESET, bus_07cbf505_);
input		CLK;
input		RESET;
output		bus_07cbf505_;
reg		kicker_1=1'h0;
wire		bus_3b0a4681_;
reg		kicker_2=1'h0;
wire		bus_59f4e2c3_;
reg		kicker_res=1'h0;
wire		bus_0476689f_;
wire		bus_4246d8a4_;
always @(posedge CLK)
begin
kicker_1<=bus_3b0a4681_;
end
assign bus_3b0a4681_=~RESET;
always @(posedge CLK)
begin
kicker_2<=bus_0476689f_;
end
assign bus_59f4e2c3_=kicker_1&bus_3b0a4681_&bus_4246d8a4_;
always @(posedge CLK)
begin
kicker_res<=bus_59f4e2c3_;
end
assign bus_07cbf505_=kicker_res;
assign bus_0476689f_=bus_3b0a4681_&kicker_1;
assign bus_4246d8a4_=~kicker_2;
endmodule



module LL2_iunzip_streamEndFun1(CLK, RESET, GO, port_27264123_, port_2c516464_, port_5613faef_, port_20d55f53_, port_0a0c52a4_, RESULT, RESULT_u950, RESULT_u951, RESULT_u952, RESULT_u953, RESULT_u954, RESULT_u955, RESULT_u956, RESULT_u957, RESULT_u958, RESULT_u959, RESULT_u960, RESULT_u961, RESULT_u962, DONE);
input		CLK;
input		RESET;
input		GO;
input		port_27264123_;
input		port_2c516464_;
input	[15:0]	port_5613faef_;
input		port_20d55f53_;
input	[15:0]	port_0a0c52a4_;
output		RESULT;
output		RESULT_u950;
output		RESULT_u951;
output	[31:0]	RESULT_u952;
output	[2:0]	RESULT_u953;
output		RESULT_u954;
output	[31:0]	RESULT_u955;
output	[2:0]	RESULT_u956;
output	[15:0]	RESULT_u957;
output	[15:0]	RESULT_u958;
output		RESULT_u959;
output		RESULT_u960;
output	[15:0]	RESULT_u961;
output	[15:0]	RESULT_u962;
output		DONE;
wire	[31:0]	add;
wire		and_u1582_u0;
wire	[8:0]	subtract;
wire		greaterThanEqualTo;
wire signed	[8:0]	greaterThanEqualTo_b_signed;
wire signed	[8:0]	greaterThanEqualTo_a_signed;
wire		and_u1583_u0;
wire		not_u308_u0;
wire		and_u1584_u0;
wire	[8:0]	subtract_u12;
wire		and_u1585_u0;
wire	[8:0]	mux_u146;
wire		and_u1586_u0;
wire	[31:0]	add_u50;
wire		and_u1587_u0;
wire		and_u1589_u0;
wire	[16:0]	add_u51;
wire	[15:0]	subtract_u13;
wire		simplePinWrite;
wire	[15:0]	simplePinWrite_u272;
wire	[15:0]	simplePinWrite_u273;
wire		simplePinWrite_u274;
wire	[15:0]	simplePinWrite_u275;
wire	[15:0]	simplePinWrite_u276;
reg		reg_249d2e91_u0=1'h0;
reg	[15:0]	syncEnable_u140=16'h0;
wire	[31:0]	mux_u147_u0;
wire		or_u430_u0;
reg	[31:0]	syncEnable_u141_u0=32'h0;
reg	[31:0]	syncEnable_u142_u0=32'h0;
reg	[15:0]	syncEnable_u143_u0=16'h0;
reg		reg_535f0a11_u0=1'h0;
assign add={31'b0, port_27264123_}+32'h0;
assign and_u1582_u0=reg_535f0a11_u0&port_2c516464_;
assign subtract={8'b0, port_27264123_}-9'h1;
assign greaterThanEqualTo_a_signed={subtract[2], subtract[2], subtract[2], subtract[2], subtract[2], subtract[2], subtract[2:0]};
assign greaterThanEqualTo_b_signed=9'h0;
assign greaterThanEqualTo=greaterThanEqualTo_a_signed>=greaterThanEqualTo_b_signed;
assign and_u1583_u0=GO&not_u308_u0;
assign not_u308_u0=~greaterThanEqualTo;
assign and_u1584_u0=GO&greaterThanEqualTo;
assign subtract_u12={8'b0, port_27264123_}-9'h1;
assign and_u1585_u0=and_u1583_u0&GO;
assign mux_u146=(and_u1585_u0)?9'h2:{subtract_u12[2], subtract_u12[2], subtract_u12[2], subtract_u12[2], subtract_u12[2], subtract_u12[2], subtract_u12[2:0]};
assign and_u1586_u0=and_u1584_u0&GO;
assign add_u50={mux_u146[2], mux_u146[2], mux_u146[2], mux_u146[2], mux_u146[2], mux_u146[2], mux_u146[2], mux_u146[2], mux_u146[2], mux_u146[2], mux_u146[2], mux_u146[2], mux_u146[2], mux_u146[2], mux_u146[2], mux_u146[2], mux_u146[2], mux_u146[2], mux_u146[2], mux_u146[2], mux_u146[2], mux_u146[2], mux_u146[2], mux_u146[2], mux_u146[2], mux_u146[2], mux_u146[2], mux_u146[2], mux_u146[2], mux_u146[2:0]}+32'h0;
assign and_u1587_u0=reg_535f0a11_u0&port_20d55f53_;
assign and_u1589_u0=reg_249d2e91_u0&port_2c516464_;
assign add_u51={syncEnable_u143_u0[15], syncEnable_u143_u0}+{port_5613faef_[15], port_5613faef_};
assign subtract_u13=syncEnable_u140-add_u51[16:1];
assign simplePinWrite=reg_249d2e91_u0&{1{reg_249d2e91_u0}};
assign simplePinWrite_u272=16'h1&{16{1'h1}};
assign simplePinWrite_u273=subtract_u13&{16{reg_249d2e91_u0}};
assign simplePinWrite_u274=reg_249d2e91_u0&{1{reg_249d2e91_u0}};
assign simplePinWrite_u275=16'h1&{16{1'h1}};
assign simplePinWrite_u276=subtract_u13&{16{reg_249d2e91_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_249d2e91_u0<=1'h0;
else reg_249d2e91_u0<=reg_535f0a11_u0;
end
always @(posedge CLK)
begin
if (reg_535f0a11_u0)
syncEnable_u140<=port_5613faef_;
end
assign mux_u147_u0=(reg_535f0a11_u0)?syncEnable_u141_u0:32'h0;
assign or_u430_u0=reg_535f0a11_u0|reg_249d2e91_u0;
always @(posedge CLK)
begin
if (GO)
syncEnable_u141_u0<={add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2:0]};
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u142_u0<=add_u50;
end
always @(posedge CLK)
begin
if (reg_535f0a11_u0)
syncEnable_u143_u0<=port_0a0c52a4_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_535f0a11_u0<=1'h0;
else reg_535f0a11_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u950=1'h0;
assign RESULT_u951=or_u430_u0;
assign RESULT_u952=mux_u147_u0;
assign RESULT_u953=3'h1;
assign RESULT_u954=reg_535f0a11_u0;
assign RESULT_u955=syncEnable_u142_u0;
assign RESULT_u956=3'h1;
assign RESULT_u957=simplePinWrite_u275;
assign RESULT_u958=simplePinWrite_u273;
assign RESULT_u959=simplePinWrite;
assign RESULT_u960=simplePinWrite_u274;
assign RESULT_u961=simplePinWrite_u272;
assign RESULT_u962=simplePinWrite_u276;
assign DONE=reg_249d2e91_u0;
endmodule



module LL2_iunzip_endianswapper_1443ed66_(endianswapper_1443ed66_in, endianswapper_1443ed66_out);
input	[31:0]	endianswapper_1443ed66_in;
output	[31:0]	endianswapper_1443ed66_out;
assign endianswapper_1443ed66_out=endianswapper_1443ed66_in;
endmodule



module LL2_iunzip_endianswapper_13a07ccf_(endianswapper_13a07ccf_in, endianswapper_13a07ccf_out);
input	[31:0]	endianswapper_13a07ccf_in;
output	[31:0]	endianswapper_13a07ccf_out;
assign endianswapper_13a07ccf_out=endianswapper_13a07ccf_in;
endmodule



module LL2_iunzip_stateVar_In1TokenIndex(bus_221c1ac8_, bus_4e95ce1d_, bus_119618fb_, bus_339b4303_, bus_32c38fb2_);
input		bus_221c1ac8_;
input		bus_4e95ce1d_;
input		bus_119618fb_;
input	[31:0]	bus_339b4303_;
output	[31:0]	bus_32c38fb2_;
wire	[31:0]	endianswapper_1443ed66_out;
reg	[31:0]	stateVar_In1TokenIndex_u2=32'h0;
wire	[31:0]	endianswapper_13a07ccf_out;
LL2_iunzip_endianswapper_1443ed66_ LL2_iunzip_endianswapper_1443ed66__1(.endianswapper_1443ed66_in(stateVar_In1TokenIndex_u2), 
  .endianswapper_1443ed66_out(endianswapper_1443ed66_out));
assign bus_32c38fb2_=endianswapper_1443ed66_out;
always @(posedge bus_221c1ac8_ or posedge bus_4e95ce1d_)
begin
if (bus_4e95ce1d_)
stateVar_In1TokenIndex_u2<=32'h0;
else if (bus_119618fb_)
stateVar_In1TokenIndex_u2<=endianswapper_13a07ccf_out;
end
LL2_iunzip_endianswapper_13a07ccf_ LL2_iunzip_endianswapper_13a07ccf__1(.endianswapper_13a07ccf_in(bus_339b4303_), 
  .endianswapper_13a07ccf_out(endianswapper_13a07ccf_out));
endmodule



module LL2_iunzip_endianswapper_4f1114ca_(endianswapper_4f1114ca_in, endianswapper_4f1114ca_out);
input	[31:0]	endianswapper_4f1114ca_in;
output	[31:0]	endianswapper_4f1114ca_out;
assign endianswapper_4f1114ca_out=endianswapper_4f1114ca_in;
endmodule



module LL2_iunzip_endianswapper_026a5845_(endianswapper_026a5845_in, endianswapper_026a5845_out);
input	[31:0]	endianswapper_026a5845_in;
output	[31:0]	endianswapper_026a5845_out;
assign endianswapper_026a5845_out={endianswapper_026a5845_in[31:2], 1'b1, endianswapper_026a5845_in[0]};
endmodule



module LL2_iunzip_stateVar_In1MaxTokenIndex(bus_54c26aa4_, bus_19793f6e_, bus_299324f7_, bus_3e112cd2_, bus_0e817a69_);
input		bus_54c26aa4_;
input		bus_19793f6e_;
input		bus_299324f7_;
input	[31:0]	bus_3e112cd2_;
output	[31:0]	bus_0e817a69_;
reg	[31:0]	stateVar_In1MaxTokenIndex_u2=32'h0;
wire	[31:0]	endianswapper_4f1114ca_out;
wire	[31:0]	endianswapper_026a5845_out;
always @(posedge bus_54c26aa4_ or posedge bus_19793f6e_)
begin
if (bus_19793f6e_)
stateVar_In1MaxTokenIndex_u2<=32'h0;
else if (bus_299324f7_)
stateVar_In1MaxTokenIndex_u2<={endianswapper_026a5845_out[31:2], 1'b1, endianswapper_026a5845_out[0]};
end
assign bus_0e817a69_=endianswapper_4f1114ca_out;
LL2_iunzip_endianswapper_4f1114ca_ LL2_iunzip_endianswapper_4f1114ca__1(.endianswapper_4f1114ca_in(stateVar_In1MaxTokenIndex_u2), 
  .endianswapper_4f1114ca_out(endianswapper_4f1114ca_out));
LL2_iunzip_endianswapper_026a5845_ LL2_iunzip_endianswapper_026a5845__1(.endianswapper_026a5845_in({bus_3e112cd2_[31:2], 1'b0, bus_3e112cd2_[0]}), 
  .endianswapper_026a5845_out(endianswapper_026a5845_out));
endmodule



module LL2_iunzip_endianswapper_78e9c6b8_(endianswapper_78e9c6b8_in, endianswapper_78e9c6b8_out);
input	[1:0]	endianswapper_78e9c6b8_in;
output	[1:0]	endianswapper_78e9c6b8_out;
assign endianswapper_78e9c6b8_out=endianswapper_78e9c6b8_in;
endmodule



module LL2_iunzip_endianswapper_0142cc2e_(endianswapper_0142cc2e_in, endianswapper_0142cc2e_out);
input	[1:0]	endianswapper_0142cc2e_in;
output	[1:0]	endianswapper_0142cc2e_out;
assign endianswapper_0142cc2e_out=endianswapper_0142cc2e_in;
endmodule



module LL2_iunzip_stateVar_fsmState_LL2_iunzip(bus_2d067e63_, bus_38ab1e34_, bus_3d48ec63_, bus_43199831_, bus_3c983ce7_);
input		bus_2d067e63_;
input		bus_38ab1e34_;
input		bus_3d48ec63_;
input	[1:0]	bus_43199831_;
output	[1:0]	bus_3c983ce7_;
wire	[1:0]	endianswapper_78e9c6b8_out;
reg	[1:0]	stateVar_fsmState_LL2_iunzip_u0=2'h0;
wire	[1:0]	endianswapper_0142cc2e_out;
LL2_iunzip_endianswapper_78e9c6b8_ LL2_iunzip_endianswapper_78e9c6b8__1(.endianswapper_78e9c6b8_in(stateVar_fsmState_LL2_iunzip_u0), 
  .endianswapper_78e9c6b8_out(endianswapper_78e9c6b8_out));
assign bus_3c983ce7_=endianswapper_78e9c6b8_out;
always @(posedge bus_2d067e63_ or posedge bus_38ab1e34_)
begin
if (bus_38ab1e34_)
stateVar_fsmState_LL2_iunzip_u0<=2'h0;
else if (bus_3d48ec63_)
stateVar_fsmState_LL2_iunzip_u0<=endianswapper_0142cc2e_out;
end
LL2_iunzip_endianswapper_0142cc2e_ LL2_iunzip_endianswapper_0142cc2e__1(.endianswapper_0142cc2e_in(bus_43199831_), 
  .endianswapper_0142cc2e_out(endianswapper_0142cc2e_out));
endmodule



module LL2_iunzip_endianswapper_49421f9e_(endianswapper_49421f9e_in, endianswapper_49421f9e_out);
input	[31:0]	endianswapper_49421f9e_in;
output	[31:0]	endianswapper_49421f9e_out;
assign endianswapper_49421f9e_out=endianswapper_49421f9e_in;
endmodule



module LL2_iunzip_endianswapper_6257f44a_(endianswapper_6257f44a_in, endianswapper_6257f44a_out);
input	[31:0]	endianswapper_6257f44a_in;
output	[31:0]	endianswapper_6257f44a_out;
assign endianswapper_6257f44a_out=endianswapper_6257f44a_in;
endmodule



module LL2_iunzip_stateVar_consumed(bus_416e1293_, bus_12087713_, bus_191cf97c_, bus_79b6c0b0_, bus_3df41d15_, bus_6619539b_, bus_5630e916_, bus_7ed235d5_, bus_13fc03a5_);
input		bus_416e1293_;
input		bus_12087713_;
input		bus_191cf97c_;
input	[31:0]	bus_79b6c0b0_;
input		bus_3df41d15_;
input	[31:0]	bus_6619539b_;
input		bus_5630e916_;
input	[31:0]	bus_7ed235d5_;
output	[31:0]	bus_13fc03a5_;
wire		or_4baa0649_u0;
wire	[31:0]	mux_1ff9c9e2_u0;
wire	[31:0]	endianswapper_49421f9e_out;
wire	[31:0]	endianswapper_6257f44a_out;
reg	[31:0]	stateVar_consumed_u4=32'h0;
assign or_4baa0649_u0=bus_191cf97c_|bus_3df41d15_|bus_5630e916_;
assign bus_13fc03a5_=endianswapper_49421f9e_out;
assign mux_1ff9c9e2_u0=({32{bus_191cf97c_}}&bus_79b6c0b0_)|({32{bus_3df41d15_}}&bus_6619539b_)|({32{bus_5630e916_}}&bus_7ed235d5_);
LL2_iunzip_endianswapper_49421f9e_ LL2_iunzip_endianswapper_49421f9e__1(.endianswapper_49421f9e_in(stateVar_consumed_u4), 
  .endianswapper_49421f9e_out(endianswapper_49421f9e_out));
LL2_iunzip_endianswapper_6257f44a_ LL2_iunzip_endianswapper_6257f44a__1(.endianswapper_6257f44a_in(mux_1ff9c9e2_u0), 
  .endianswapper_6257f44a_out(endianswapper_6257f44a_out));
always @(posedge bus_416e1293_ or posedge bus_12087713_)
begin
if (bus_12087713_)
stateVar_consumed_u4<=32'h0;
else if (or_4baa0649_u0)
stateVar_consumed_u4<=endianswapper_6257f44a_out;
end
endmodule



module LL2_iunzip_streamEndFun2(CLK, RESET, GO, port_2a8e19bd_, port_377c7b5e_, port_3606eb83_, port_1d8d2ce2_, port_2bdba753_, RESULT, RESULT_u963, RESULT_u964, RESULT_u965, RESULT_u966, RESULT_u967, RESULT_u968, RESULT_u969, RESULT_u970, RESULT_u971, RESULT_u972, RESULT_u973, RESULT_u974, RESULT_u975, DONE);
input		CLK;
input		RESET;
input		GO;
input		port_2a8e19bd_;
input		port_377c7b5e_;
input	[15:0]	port_3606eb83_;
input		port_1d8d2ce2_;
input	[15:0]	port_2bdba753_;
output		RESULT;
output		RESULT_u963;
output		RESULT_u964;
output	[31:0]	RESULT_u965;
output	[2:0]	RESULT_u966;
output		RESULT_u967;
output	[31:0]	RESULT_u968;
output	[2:0]	RESULT_u969;
output	[15:0]	RESULT_u970;
output	[15:0]	RESULT_u971;
output		RESULT_u972;
output		RESULT_u973;
output	[15:0]	RESULT_u974;
output	[15:0]	RESULT_u975;
output		DONE;
wire	[31:0]	add;
wire		and_u1591_u0;
wire	[8:0]	subtract;
wire signed	[8:0]	greaterThanEqualTo_a_signed;
wire		greaterThanEqualTo;
wire signed	[8:0]	greaterThanEqualTo_b_signed;
wire		not_u309_u0;
wire		and_u1592_u0;
wire		and_u1593_u0;
wire	[8:0]	subtract_u14;
wire		and_u1594_u0;
wire		and_u1595_u0;
wire	[8:0]	mux_u148;
wire	[31:0]	add_u52;
wire		and_u1596_u0;
wire		and_u1598_u0;
wire	[16:0]	add_u53;
wire	[15:0]	add_u54;
wire		simplePinWrite;
wire	[15:0]	simplePinWrite_u277;
wire	[15:0]	simplePinWrite_u278;
wire	[15:0]	simplePinWrite_u279;
wire		simplePinWrite_u280;
wire	[15:0]	simplePinWrite_u281;
reg		reg_62440bcd_u0=1'h0;
reg	[15:0]	syncEnable_u144=16'h0;
reg	[31:0]	syncEnable_u145_u0=32'h0;
reg		reg_245abd9f_u0=1'h0;
reg	[15:0]	syncEnable_u146_u0=16'h0;
reg	[31:0]	syncEnable_u147_u0=32'h0;
wire	[31:0]	mux_u149_u0;
wire		or_u431_u0;
assign add={31'b0, port_2a8e19bd_}+32'h0;
assign and_u1591_u0=reg_245abd9f_u0&port_377c7b5e_;
assign subtract={8'b0, port_2a8e19bd_}-9'h1;
assign greaterThanEqualTo_a_signed={subtract[2], subtract[2], subtract[2], subtract[2], subtract[2], subtract[2], subtract[2:0]};
assign greaterThanEqualTo_b_signed=9'h0;
assign greaterThanEqualTo=greaterThanEqualTo_a_signed>=greaterThanEqualTo_b_signed;
assign not_u309_u0=~greaterThanEqualTo;
assign and_u1592_u0=GO&greaterThanEqualTo;
assign and_u1593_u0=GO&not_u309_u0;
assign subtract_u14={8'b0, port_2a8e19bd_}-9'h1;
assign and_u1594_u0=and_u1592_u0&GO;
assign and_u1595_u0=and_u1593_u0&GO;
assign mux_u148=(and_u1594_u0)?{subtract_u14[2], subtract_u14[2], subtract_u14[2], subtract_u14[2], subtract_u14[2], subtract_u14[2], subtract_u14[2:0]}:9'h2;
assign add_u52={mux_u148[2], mux_u148[2], mux_u148[2], mux_u148[2], mux_u148[2], mux_u148[2], mux_u148[2], mux_u148[2], mux_u148[2], mux_u148[2], mux_u148[2], mux_u148[2], mux_u148[2], mux_u148[2], mux_u148[2], mux_u148[2], mux_u148[2], mux_u148[2], mux_u148[2], mux_u148[2], mux_u148[2], mux_u148[2], mux_u148[2], mux_u148[2], mux_u148[2], mux_u148[2], mux_u148[2], mux_u148[2], mux_u148[2], mux_u148[2:0]}+32'h0;
assign and_u1596_u0=reg_245abd9f_u0&port_1d8d2ce2_;
assign and_u1598_u0=reg_62440bcd_u0&port_377c7b5e_;
assign add_u53={syncEnable_u146_u0[15], syncEnable_u146_u0}+{port_3606eb83_[15], port_3606eb83_};
assign add_u54=syncEnable_u144+{add_u53[16], add_u53[16:2]};
assign simplePinWrite=reg_62440bcd_u0&{1{reg_62440bcd_u0}};
assign simplePinWrite_u277=add_u54&{16{reg_62440bcd_u0}};
assign simplePinWrite_u278=16'h1&{16{1'h1}};
assign simplePinWrite_u279=16'h1&{16{1'h1}};
assign simplePinWrite_u280=reg_62440bcd_u0&{1{reg_62440bcd_u0}};
assign simplePinWrite_u281=add_u54&{16{reg_62440bcd_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_62440bcd_u0<=1'h0;
else reg_62440bcd_u0<=reg_245abd9f_u0;
end
always @(posedge CLK)
begin
if (reg_245abd9f_u0)
syncEnable_u144<=port_3606eb83_;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u145_u0<=add_u52;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_245abd9f_u0<=1'h0;
else reg_245abd9f_u0<=GO;
end
always @(posedge CLK)
begin
if (reg_245abd9f_u0)
syncEnable_u146_u0<=port_2bdba753_;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u147_u0<={add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2:0]};
end
assign mux_u149_u0=(reg_245abd9f_u0)?syncEnable_u147_u0:32'h0;
assign or_u431_u0=reg_245abd9f_u0|reg_62440bcd_u0;
assign RESULT=GO;
assign RESULT_u963=1'h0;
assign RESULT_u964=or_u431_u0;
assign RESULT_u965=mux_u149_u0;
assign RESULT_u966=3'h1;
assign RESULT_u967=reg_245abd9f_u0;
assign RESULT_u968=syncEnable_u145_u0;
assign RESULT_u969=3'h1;
assign RESULT_u970=simplePinWrite_u279;
assign RESULT_u971=simplePinWrite_u277;
assign RESULT_u972=simplePinWrite;
assign RESULT_u973=simplePinWrite_u280;
assign RESULT_u974=simplePinWrite_u278;
assign RESULT_u975=simplePinWrite_u281;
assign DONE=reg_62440bcd_u0;
endmodule



module LL2_iunzip_endianswapper_1ba7c737_(endianswapper_1ba7c737_in, endianswapper_1ba7c737_out);
input	[1:0]	endianswapper_1ba7c737_in;
output	[1:0]	endianswapper_1ba7c737_out;
assign endianswapper_1ba7c737_out=endianswapper_1ba7c737_in;
endmodule



module LL2_iunzip_endianswapper_539905b2_(endianswapper_539905b2_in, endianswapper_539905b2_out);
input	[1:0]	endianswapper_539905b2_in;
output	[1:0]	endianswapper_539905b2_out;
assign endianswapper_539905b2_out=endianswapper_539905b2_in;
endmodule



module LL2_iunzip_stateVar_fsmOldState_LL2_iunzip(bus_3b581e33_, bus_52d5710c_, bus_4ec3c878_, bus_4cb5a4aa_, bus_3078af4b_);
input		bus_3b581e33_;
input		bus_52d5710c_;
input		bus_4ec3c878_;
input	[1:0]	bus_4cb5a4aa_;
output	[1:0]	bus_3078af4b_;
wire	[1:0]	endianswapper_1ba7c737_out;
reg	[1:0]	stateVar_fsmOldState_LL2_iunzip_u0=2'h0;
wire	[1:0]	endianswapper_539905b2_out;
LL2_iunzip_endianswapper_1ba7c737_ LL2_iunzip_endianswapper_1ba7c737__1(.endianswapper_1ba7c737_in(bus_4cb5a4aa_), 
  .endianswapper_1ba7c737_out(endianswapper_1ba7c737_out));
always @(posedge bus_3b581e33_ or posedge bus_52d5710c_)
begin
if (bus_52d5710c_)
stateVar_fsmOldState_LL2_iunzip_u0<=2'h0;
else if (bus_4ec3c878_)
stateVar_fsmOldState_LL2_iunzip_u0<=endianswapper_1ba7c737_out;
end
LL2_iunzip_endianswapper_539905b2_ LL2_iunzip_endianswapper_539905b2__1(.endianswapper_539905b2_in(stateVar_fsmOldState_LL2_iunzip_u0), 
  .endianswapper_539905b2_out(endianswapper_539905b2_out));
assign bus_3078af4b_=endianswapper_539905b2_out;
endmodule



module LL2_iunzip_streamFun2(CLK, RESET, GO, port_5fca059d_, port_581d88d1_, port_79fe3347_, port_3b68465d_, port_7396b25e_, port_33e93e76_, port_4ccd3ea3_, port_2d7037ba_, RESULT, RESULT_u976, RESULT_u977, RESULT_u978, RESULT_u979, RESULT_u980, RESULT_u981, RESULT_u982, RESULT_u983, RESULT_u984, RESULT_u985, RESULT_u986, RESULT_u987, RESULT_u988, RESULT_u989, RESULT_u990, RESULT_u991, RESULT_u992, DONE);
input		CLK;
input		RESET;
input		GO;
input		port_5fca059d_;
input	[31:0]	port_581d88d1_;
input		port_79fe3347_;
input	[15:0]	port_3b68465d_;
input		port_7396b25e_;
input	[15:0]	port_33e93e76_;
input		port_4ccd3ea3_;
input	[15:0]	port_2d7037ba_;
output		RESULT;
output		RESULT_u976;
output		RESULT_u977;
output	[31:0]	RESULT_u978;
output		RESULT_u979;
output	[31:0]	RESULT_u980;
output	[2:0]	RESULT_u981;
output		RESULT_u982;
output	[31:0]	RESULT_u983;
output	[2:0]	RESULT_u984;
output		RESULT_u985;
output	[31:0]	RESULT_u986;
output	[15:0]	RESULT_u987;
output	[2:0]	RESULT_u988;
output	[15:0]	RESULT_u989;
output		RESULT_u990;
output		RESULT_u991;
output	[15:0]	RESULT_u992;
output		DONE;
wire		simplePinWrite;
reg		reg_76dec11f_u0=1'h0;
wire		or_u432_u0;
wire		and_u1601_u0;
wire	[31:0]	add;
wire		and_u1602_u0;
wire	[8:0]	subtract;
wire signed	[8:0]	greaterThanEqualTo_b_signed;
wire signed	[8:0]	greaterThanEqualTo_a_signed;
wire		greaterThanEqualTo;
wire		not_u310_u0;
wire		and_u1603_u0;
wire		and_u1604_u0;
wire	[8:0]	subtract_u15;
wire		and_u1605_u0;
wire		and_u1606_u0;
wire	[8:0]	mux_u150;
wire	[31:0]	add_u55;
wire		and_u1607_u0;
wire		and_u1609_u0;
wire	[16:0]	add_u56;
wire	[15:0]	add_u57;
wire	[31:0]	add_u58;
wire		simplePinWrite_u282;
wire	[15:0]	simplePinWrite_u283;
wire	[15:0]	simplePinWrite_u284;
reg	[31:0]	syncEnable_u148=32'h0;
reg	[15:0]	syncEnable_u149_u0=16'h0;
reg		reg_7a8b9ad9_u0=1'h0;
wire		or_u433_u0;
wire	[31:0]	mux_u151_u0;
reg		reg_7a8b9ad9_result_delayed_u0=1'h0;
reg	[31:0]	syncEnable_u150_u0=32'h0;
wire	[31:0]	mux_u152_u0;
reg	[15:0]	syncEnable_u151_u0=16'h0;
reg	[15:0]	syncEnable_u152_u0=16'h0;
reg		reg_7a8b9ad9_result_delayed_result_delayed_u0=1'h0;
assign simplePinWrite=GO&{1{GO}};
always @(posedge CLK or posedge reg_7a8b9ad9_u0 or posedge or_u432_u0)
begin
if (or_u432_u0)
reg_76dec11f_u0<=1'h0;
else if (reg_7a8b9ad9_u0)
reg_76dec11f_u0<=1'h1;
else reg_76dec11f_u0<=reg_76dec11f_u0;
end
assign or_u432_u0=and_u1601_u0|RESET;
assign and_u1601_u0=reg_76dec11f_u0&port_4ccd3ea3_;
assign add={31'b0, port_5fca059d_}+32'h0;
assign and_u1602_u0=reg_7a8b9ad9_result_delayed_u0&port_79fe3347_;
assign subtract={8'b0, port_5fca059d_}-9'h1;
assign greaterThanEqualTo_a_signed={subtract[2], subtract[2], subtract[2], subtract[2], subtract[2], subtract[2], subtract[2:0]};
assign greaterThanEqualTo_b_signed=9'h0;
assign greaterThanEqualTo=greaterThanEqualTo_a_signed>=greaterThanEqualTo_b_signed;
assign not_u310_u0=~greaterThanEqualTo;
assign and_u1603_u0=GO&greaterThanEqualTo;
assign and_u1604_u0=GO&not_u310_u0;
assign subtract_u15={8'b0, port_5fca059d_}-9'h1;
assign and_u1605_u0=and_u1603_u0&GO;
assign and_u1606_u0=and_u1604_u0&GO;
assign mux_u150=(and_u1606_u0)?9'h2:{subtract_u15[2], subtract_u15[2], subtract_u15[2], subtract_u15[2], subtract_u15[2], subtract_u15[2], subtract_u15[2:0]};
assign add_u55={mux_u150[2], mux_u150[2], mux_u150[2], mux_u150[2], mux_u150[2], mux_u150[2], mux_u150[2], mux_u150[2], mux_u150[2], mux_u150[2], mux_u150[2], mux_u150[2], mux_u150[2], mux_u150[2], mux_u150[2], mux_u150[2], mux_u150[2], mux_u150[2], mux_u150[2], mux_u150[2], mux_u150[2], mux_u150[2], mux_u150[2], mux_u150[2], mux_u150[2], mux_u150[2], mux_u150[2], mux_u150[2], mux_u150[2], mux_u150[2:0]}+32'h0;
assign and_u1607_u0=reg_7a8b9ad9_result_delayed_u0&port_4ccd3ea3_;
assign and_u1609_u0=reg_7a8b9ad9_result_delayed_result_delayed_u0&port_79fe3347_;
assign add_u56={syncEnable_u151_u0[15], syncEnable_u151_u0}+{port_3b68465d_[15], port_3b68465d_};
assign add_u57=syncEnable_u149_u0+{add_u56[16], add_u56[16:2]};
assign add_u58=port_581d88d1_+32'h1;
assign simplePinWrite_u282=reg_7a8b9ad9_result_delayed_result_delayed_u0&{1{reg_7a8b9ad9_result_delayed_result_delayed_u0}};
assign simplePinWrite_u283=add_u57&{16{reg_7a8b9ad9_result_delayed_result_delayed_u0}};
assign simplePinWrite_u284=16'h1&{16{1'h1}};
always @(posedge CLK)
begin
if (GO)
syncEnable_u148<={add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2:0]};
end
always @(posedge CLK)
begin
if (reg_7a8b9ad9_result_delayed_u0)
syncEnable_u149_u0<=port_3b68465d_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a8b9ad9_u0<=1'h0;
else reg_7a8b9ad9_u0<=GO;
end
assign or_u433_u0=reg_7a8b9ad9_result_delayed_u0|reg_7a8b9ad9_result_delayed_result_delayed_u0;
assign mux_u151_u0=(reg_7a8b9ad9_result_delayed_u0)?syncEnable_u148:32'h0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a8b9ad9_result_delayed_u0<=1'h0;
else reg_7a8b9ad9_result_delayed_u0<=reg_7a8b9ad9_u0;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u150_u0<=add_u55;
end
assign mux_u152_u0=(reg_7a8b9ad9_u0)?32'h0:syncEnable_u150_u0;
always @(posedge CLK)
begin
if (reg_7a8b9ad9_result_delayed_u0)
syncEnable_u151_u0<=port_33e93e76_;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u152_u0<=port_2d7037ba_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a8b9ad9_result_delayed_result_delayed_u0<=1'h0;
else reg_7a8b9ad9_result_delayed_result_delayed_u0<=reg_7a8b9ad9_result_delayed_u0;
end
assign RESULT=GO;
assign RESULT_u976=1'h0;
assign RESULT_u977=GO;
assign RESULT_u978=add_u58;
assign RESULT_u979=or_u433_u0;
assign RESULT_u980=mux_u151_u0;
assign RESULT_u981=3'h1;
assign RESULT_u982=reg_7a8b9ad9_result_delayed_u0;
assign RESULT_u983=mux_u152_u0;
assign RESULT_u984=3'h1;
assign RESULT_u985=reg_7a8b9ad9_u0;
assign RESULT_u986=mux_u152_u0;
assign RESULT_u987=syncEnable_u152_u0;
assign RESULT_u988=3'h1;
assign RESULT_u989=simplePinWrite_u284;
assign RESULT_u990=simplePinWrite_u282;
assign RESULT_u991=simplePinWrite;
assign RESULT_u992=simplePinWrite_u283;
assign DONE=reg_7a8b9ad9_result_delayed_result_delayed_u0;
endmodule



module LL2_iunzip_simplememoryreferee_15caad00_(bus_16cdabb7_, bus_0de57dc4_, bus_7b32a18c_, bus_247edfb6_, bus_229405ff_, bus_5a473665_, bus_36b4444a_, bus_005f3f40_, bus_1d7ad841_, bus_36f7a4bd_, bus_6d1b31d9_, bus_7046b040_, bus_6715655d_, bus_1d3acc5f_);
input		bus_16cdabb7_;
input		bus_0de57dc4_;
input		bus_7b32a18c_;
input	[15:0]	bus_247edfb6_;
input		bus_229405ff_;
input	[31:0]	bus_5a473665_;
input	[2:0]	bus_36b4444a_;
output	[15:0]	bus_005f3f40_;
output	[31:0]	bus_1d7ad841_;
output		bus_36f7a4bd_;
output		bus_6d1b31d9_;
output	[2:0]	bus_7046b040_;
output	[15:0]	bus_6715655d_;
output		bus_1d3acc5f_;
assign bus_005f3f40_=16'h0;
assign bus_1d7ad841_=32'h1;
assign bus_36f7a4bd_=1'h0;
assign bus_6d1b31d9_=bus_229405ff_;
assign bus_7046b040_=3'h1;
assign bus_6715655d_=bus_247edfb6_;
assign bus_1d3acc5f_=bus_7b32a18c_;
endmodule



module LL2_iunzip_forge_memory_2x16_15(CLK, ENA, WEA, DINA, ENB, ADDRA, ADDRB, DOUTA, DOUTB, DONEA, DONEB);
input		CLK;
input		ENA;
input		WEA;
input	[15:0]	DINA;
input		ENB;
input	[31:0]	ADDRA;
input	[31:0]	ADDRB;
output	[15:0]	DOUTA;
output	[15:0]	DOUTB;
output		DONEA;
output		DONEB;
wire		wea_0;
wire	[15:0]	pre_douta_0;
wire	[15:0]	pre_doutb_0;
reg		wea_done;
reg		rea_done;
reg	[15:0]	mux_outa;
reg	[15:0]	mux_outb;
assign wea_0=WEA;
always @(posedge CLK)
begin
wea_done<=WEA;
end
assign DONEA=rea_done|wea_done;
always @(posedge CLK)
begin
end
assign DONEB=ENB;
always @(pre_douta_0)
begin
mux_outa<=pre_douta_0;
end
assign DOUTA=mux_outa;
always @(pre_doutb_0)
begin
mux_outb<=pre_doutb_0;
end
assign DOUTB=mux_outb;
// Memory array element: COL: 0, ROW: 0
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_80(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[0]), .SPO(pre_douta_0[0]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[0]));
// Memory array element: COL: 0, ROW: 1
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_81(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[1]), .SPO(pre_douta_0[1]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[1]));
// Memory array element: COL: 0, ROW: 2
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_82(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[2]), .SPO(pre_douta_0[2]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[2]));
// Memory array element: COL: 0, ROW: 3
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_83(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[3]), .SPO(pre_douta_0[3]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[3]));
// Memory array element: COL: 0, ROW: 4
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_84(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[4]), .SPO(pre_douta_0[4]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[4]));
// Memory array element: COL: 0, ROW: 5
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_85(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[5]), .SPO(pre_douta_0[5]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[5]));
// Memory array element: COL: 0, ROW: 6
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_86(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[6]), .SPO(pre_douta_0[6]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[6]));
// Memory array element: COL: 0, ROW: 7
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_87(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[7]), .SPO(pre_douta_0[7]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[7]));
// Memory array element: COL: 0, ROW: 8
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_88(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[8]), .SPO(pre_douta_0[8]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[8]));
// Memory array element: COL: 0, ROW: 9
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_89(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[9]), .SPO(pre_douta_0[9]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[9]));
// Memory array element: COL: 0, ROW: 10
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_90(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[10]), .SPO(pre_douta_0[10]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[10]));
// Memory array element: COL: 0, ROW: 11
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_91(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[11]), .SPO(pre_douta_0[11]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[11]));
// Memory array element: COL: 0, ROW: 12
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_92(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[12]), .SPO(pre_douta_0[12]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[12]));
// Memory array element: COL: 0, ROW: 13
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_93(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[13]), .SPO(pre_douta_0[13]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[13]));
// Memory array element: COL: 0, ROW: 14
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_94(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[14]), .SPO(pre_douta_0[14]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[14]));
// Memory array element: COL: 0, ROW: 15
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_95(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[15]), .SPO(pre_douta_0[15]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[15]));
endmodule



module LL2_iunzip_structuralmemory_0e000751_(CLK_u7, bus_457d065b_, bus_417f17f6_, bus_7399bd45_, bus_6a7bbc81_, bus_3cbe9f79_, bus_04ea2051_, bus_4640c3a2_, bus_73e3f3e7_, bus_4ce023f4_, bus_29133072_, bus_52940f8a_, bus_066c060a_, bus_0c01b8a2_);
input		CLK_u7;
input		bus_457d065b_;
input	[31:0]	bus_417f17f6_;
input	[2:0]	bus_7399bd45_;
input		bus_6a7bbc81_;
input	[31:0]	bus_3cbe9f79_;
input	[2:0]	bus_04ea2051_;
input		bus_4640c3a2_;
input		bus_73e3f3e7_;
input	[15:0]	bus_4ce023f4_;
output	[15:0]	bus_29133072_;
output		bus_52940f8a_;
output	[15:0]	bus_066c060a_;
output		bus_0c01b8a2_;
wire		or_025c90fe_u0;
wire		or_1a5243b6_u0;
wire		and_6e8649ee_u0;
reg		logicalMem_30648013_we_delay0_u0=1'h0;
wire	[15:0]	bus_0d59d088_;
wire	[15:0]	bus_4752fb7f_;
wire		not_30ac475a_u0;
assign or_025c90fe_u0=and_6e8649ee_u0|logicalMem_30648013_we_delay0_u0;
assign or_1a5243b6_u0=bus_4640c3a2_|bus_73e3f3e7_;
assign and_6e8649ee_u0=bus_4640c3a2_&not_30ac475a_u0;
always @(posedge CLK_u7 or posedge bus_457d065b_)
begin
if (bus_457d065b_)
logicalMem_30648013_we_delay0_u0<=1'h0;
else logicalMem_30648013_we_delay0_u0<=bus_73e3f3e7_;
end
assign bus_29133072_=bus_0d59d088_;
assign bus_52940f8a_=bus_6a7bbc81_;
assign bus_066c060a_=bus_4752fb7f_;
assign bus_0c01b8a2_=or_025c90fe_u0;
LL2_iunzip_forge_memory_2x16_15 LL2_iunzip_forge_memory_2x16_15_instance0(.CLK(CLK_u7), 
  .ENA(or_1a5243b6_u0), .WEA(bus_73e3f3e7_), .DINA(bus_4ce023f4_), .ADDRA(bus_3cbe9f79_), 
  .DOUTA(bus_4752fb7f_), .DONEA(), .ENB(bus_6a7bbc81_), .ADDRB(32'h1), .DOUTB(bus_0d59d088_), 
  .DONEB());
assign not_30ac475a_u0=~bus_73e3f3e7_;
endmodule



module LL2_iunzip_simplememoryreferee_06e2d637_(bus_54a19bc9_, bus_4453c8b0_, bus_567d4ed5_, bus_59677524_, bus_209bc1d3_, bus_2383042c_, bus_355229bb_, bus_765ef4b2_, bus_23a9aa5b_, bus_0d9a64c8_, bus_17a89a93_, bus_5555630d_, bus_3552a76c_, bus_57a3f872_, bus_5ee3d6e0_, bus_6483aa66_, bus_6cf5cfbb_, bus_62f7ce09_, bus_35ec3db3_, bus_27b331c3_, bus_14e11e79_, bus_6ee688b9_, bus_2284bbc7_, bus_1c9a0cac_, bus_7ca96f1c_, bus_2873baa2_, bus_7db96305_, bus_7c6d4762_, bus_79309e44_, bus_72817d63_, bus_5a3ab128_, bus_01050093_, bus_7e0b6b8d_, bus_44703396_, bus_7045541b_, bus_539df49f_, bus_5263a0f6_, bus_0e4c9451_);
input		bus_54a19bc9_;
input		bus_4453c8b0_;
input		bus_567d4ed5_;
input	[15:0]	bus_59677524_;
input		bus_209bc1d3_;
input	[15:0]	bus_2383042c_;
input	[31:0]	bus_355229bb_;
input	[2:0]	bus_765ef4b2_;
input		bus_23a9aa5b_;
input		bus_0d9a64c8_;
input	[15:0]	bus_17a89a93_;
input	[31:0]	bus_5555630d_;
input	[2:0]	bus_3552a76c_;
input		bus_57a3f872_;
input		bus_5ee3d6e0_;
input	[15:0]	bus_6483aa66_;
input	[31:0]	bus_6cf5cfbb_;
input	[2:0]	bus_62f7ce09_;
input		bus_35ec3db3_;
input	[31:0]	bus_27b331c3_;
input	[2:0]	bus_14e11e79_;
input		bus_6ee688b9_;
input	[31:0]	bus_2284bbc7_;
input	[2:0]	bus_1c9a0cac_;
output	[15:0]	bus_7ca96f1c_;
output	[31:0]	bus_2873baa2_;
output		bus_7db96305_;
output		bus_7c6d4762_;
output	[2:0]	bus_79309e44_;
output		bus_72817d63_;
output	[15:0]	bus_5a3ab128_;
output		bus_01050093_;
output	[15:0]	bus_7e0b6b8d_;
output		bus_44703396_;
output	[15:0]	bus_7045541b_;
output		bus_539df49f_;
output	[15:0]	bus_5263a0f6_;
output		bus_0e4c9451_;
wire		not_011c5d1c_u0;
wire		and_06600263_u0;
wire		not_58bc07f8_u0;
wire		not_1560b366_u0;
wire		or_5c146613_u0;
reg		done_qual_u66_u0=1'h0;
wire		and_7ae1912a_u0;
wire		or_105abf56_u0;
wire		and_45a258f2_u0;
wire		or_1f3eb56f_u0;
wire		not_54f42566_u0;
wire		or_25266f75_u0;
wire		and_2bb1b16d_u0;
reg		done_qual_u67_u0=1'h0;
wire		or_1685e566_u0;
reg		done_qual_u68_u0=1'h0;
wire		or_1db4c21e_u0;
reg		done_qual_u69_u0=1'h0;
wire		or_4db9a580_u0;
wire		and_27a7929e_u0;
wire	[15:0]	mux_1af6facc_u0;
wire	[31:0]	mux_0dc6d6bc_u0;
wire		or_504f6e33_u0;
reg		done_qual_u70_u0=1'h0;
wire		or_6107c6f9_u0;
wire		not_0dca6434_u0;
assign not_011c5d1c_u0=~bus_567d4ed5_;
assign and_06600263_u0=or_1685e566_u0&bus_567d4ed5_;
assign not_58bc07f8_u0=~bus_567d4ed5_;
assign not_1560b366_u0=~bus_567d4ed5_;
assign or_5c146613_u0=bus_209bc1d3_|done_qual_u69_u0;
always @(posedge bus_54a19bc9_)
begin
if (bus_4453c8b0_)
done_qual_u66_u0<=1'h0;
else done_qual_u66_u0<=bus_6ee688b9_;
end
assign bus_7ca96f1c_=mux_1af6facc_u0;
assign bus_2873baa2_=mux_0dc6d6bc_u0;
assign bus_7db96305_=or_504f6e33_u0;
assign bus_7c6d4762_=or_6107c6f9_u0;
assign bus_79309e44_=3'h1;
assign bus_72817d63_=and_2bb1b16d_u0;
assign bus_5a3ab128_=bus_59677524_;
assign bus_01050093_=and_45a258f2_u0;
assign bus_7e0b6b8d_=bus_59677524_;
assign bus_44703396_=and_7ae1912a_u0;
assign bus_7045541b_=bus_59677524_;
assign bus_539df49f_=and_06600263_u0;
assign bus_5263a0f6_=bus_59677524_;
assign bus_0e4c9451_=and_27a7929e_u0;
assign and_7ae1912a_u0=or_105abf56_u0&bus_567d4ed5_;
assign or_105abf56_u0=or_25266f75_u0|done_qual_u67_u0;
assign and_45a258f2_u0=or_1f3eb56f_u0&bus_567d4ed5_;
assign or_1f3eb56f_u0=or_4db9a580_u0|done_qual_u68_u0;
assign not_54f42566_u0=~bus_567d4ed5_;
assign or_25266f75_u0=bus_57a3f872_|bus_5ee3d6e0_;
assign and_2bb1b16d_u0=or_5c146613_u0&bus_567d4ed5_;
always @(posedge bus_54a19bc9_)
begin
if (bus_4453c8b0_)
done_qual_u67_u0<=1'h0;
else done_qual_u67_u0<=or_25266f75_u0;
end
assign or_1685e566_u0=bus_35ec3db3_|done_qual_u70_u0;
always @(posedge bus_54a19bc9_)
begin
if (bus_4453c8b0_)
done_qual_u68_u0<=1'h0;
else done_qual_u68_u0<=or_4db9a580_u0;
end
assign or_1db4c21e_u0=bus_6ee688b9_|done_qual_u66_u0;
always @(posedge bus_54a19bc9_)
begin
if (bus_4453c8b0_)
done_qual_u69_u0<=1'h0;
else done_qual_u69_u0<=bus_209bc1d3_;
end
assign or_4db9a580_u0=bus_23a9aa5b_|bus_0d9a64c8_;
assign and_27a7929e_u0=or_1db4c21e_u0&bus_567d4ed5_;
assign mux_1af6facc_u0=({16{bus_209bc1d3_}}&bus_2383042c_)|({16{bus_0d9a64c8_}}&bus_17a89a93_)|({16{bus_5ee3d6e0_}}&bus_6483aa66_);
assign mux_0dc6d6bc_u0=({32{bus_209bc1d3_}}&{31'b0, bus_355229bb_[0]})|({32{or_4db9a580_u0}}&bus_5555630d_)|({32{or_25266f75_u0}}&bus_6cf5cfbb_)|({32{bus_35ec3db3_}}&bus_27b331c3_)|({32{bus_6ee688b9_}}&bus_2284bbc7_);
assign or_504f6e33_u0=bus_209bc1d3_|bus_0d9a64c8_|bus_5ee3d6e0_;
always @(posedge bus_54a19bc9_)
begin
if (bus_4453c8b0_)
done_qual_u70_u0<=1'h0;
else done_qual_u70_u0<=bus_35ec3db3_;
end
assign or_6107c6f9_u0=bus_209bc1d3_|or_4db9a580_u0|or_25266f75_u0|bus_35ec3db3_|bus_6ee688b9_;
assign not_0dca6434_u0=~bus_567d4ed5_;
endmodule



module LL2_iunzip_scheduler(CLK, RESET, GO, port_44cbc7ff_, port_57df124f_, port_2710208c_, port_0dedb00e_, port_0cb02262_, port_51623660_, port_5f577b2f_, port_2d918d8b_, port_3777dab3_, port_6a679525_, port_5a872d3c_, port_1a1203bd_, port_4cbbb047_, port_59e64907_, port_5351796d_, RESULT, RESULT_u993, RESULT_u994, RESULT_u995, RESULT_u996, RESULT_u997, RESULT_u998, RESULT_u999, RESULT_u1000, RESULT_u1001, RESULT_u1002, RESULT_u1003, RESULT_u1004, RESULT_u1005, RESULT_u1006, RESULT_u1007, RESULT_u1008, RESULT_u1009, RESULT_u1010, RESULT_u1011, DONE);
input		CLK;
input		RESET;
input		GO;
input	[1:0]	port_44cbc7ff_;
input	[1:0]	port_57df124f_;
input	[31:0]	port_2710208c_;
input	[31:0]	port_0dedb00e_;
input	[31:0]	port_0cb02262_;
input		port_51623660_;
input		port_5f577b2f_;
input		port_2d918d8b_;
input		port_3777dab3_;
input		port_6a679525_;
input	[15:0]	port_5a872d3c_;
input		port_1a1203bd_;
input		port_4cbbb047_;
input		port_59e64907_;
input		port_5351796d_;
output		RESULT;
output	[1:0]	RESULT_u993;
output		RESULT_u994;
output	[1:0]	RESULT_u995;
output		RESULT_u996;
output	[31:0]	RESULT_u997;
output		RESULT_u998;
output	[31:0]	RESULT_u999;
output		RESULT_u1000;
output		RESULT_u1001;
output		RESULT_u1002;
output	[31:0]	RESULT_u1003;
output	[15:0]	RESULT_u1004;
output	[2:0]	RESULT_u1005;
output		RESULT_u1006;
output		RESULT_u1007;
output		RESULT_u1008;
output		RESULT_u1009;
output		RESULT_u1010;
output		RESULT_u1011;
output		DONE;
wire signed	[31:0]	equals_b_signed;
wire		equals;
wire signed	[31:0]	equals_a_signed;
wire signed	[31:0]	equals_u86_b_signed;
wire		equals_u86;
wire signed	[31:0]	equals_u86_a_signed;
wire		equals_u87;
wire signed	[31:0]	equals_u87_a_signed;
wire signed	[31:0]	equals_u87_b_signed;
wire signed	[31:0]	equals_u88_a_signed;
wire signed	[31:0]	equals_u88_b_signed;
wire		equals_u88;
wire		not_u311_u0;
wire		and_u1611_u0;
wire		and_u1612_u0;
wire		and_u1613_u0;
wire		not_u312_u0;
wire		and_u1614_u0;
wire		simplePinWrite;
reg		reg_077142d5_u0=1'h0;
reg		reg_077142d5_result_delayed_u0=1'h0;
wire		or_u434_u0;
reg		reg_2f7b9f51_u0=1'h0;
wire	[1:0]	mux_u153;
wire		or_u435_u0;
wire		and_u1615_u0;
wire		and_u1616_u0;
reg		and_delayed_u103=1'h0;
wire		and_u1617_u0;
wire		and_u1618_u0;
wire		or_u436_u0;
reg		and_delayed_u104_u0=1'h0;
wire signed	[31:0]	equals_u89_a_signed;
wire signed	[31:0]	equals_u89_b_signed;
wire		equals_u89;
wire		and_u1619_u0;
wire		not_u313_u0;
wire		and_u1620_u0;
wire		and_u1621_u0;
wire		and_u1622_u0;
wire		not_u314_u0;
wire		andOp;
wire		and_u1623_u0;
wire		and_u1624_u0;
wire		not_u315_u0;
wire		simplePinWrite_u285;
wire		and_u1625_u0;
wire		or_u437_u0;
reg		reg_71668bce_u0=1'h0;
reg		reg_76959641_u0=1'h0;
reg		and_delayed_u105_u0=1'h0;
wire		and_u1626_u0;
wire		and_u1627_u0;
wire		and_u1628_u0;
wire		not_u316_u0;
wire		and_u1629_u0;
wire		not_u317_u0;
wire		and_u1630_u0;
wire		simplePinWrite_u286;
wire		or_u438_u0;
reg		reg_154898a9_u0=1'h0;
wire		and_u1631_u0;
reg		and_delayed_u106_u0=1'h0;
reg		reg_7e4e1b1e_u0=1'h0;
reg		and_delayed_result_delayed_u8=1'h0;
wire		and_u1632_u0;
wire		or_u439_u0;
wire	[1:0]	mux_u154_u0;
wire		and_u1633_u0;
reg		and_delayed_u107_u0=1'h0;
wire		and_u1634_u0;
wire		or_u440_u0;
wire		and_u1635_u0;
wire		or_u441_u0;
wire	[1:0]	mux_u155_u0;
wire		and_u1636_u0;
wire		or_u442_u0;
wire		and_u1637_u0;
wire		and_u1638_u0;
wire		or_u443_u0;
reg		and_delayed_u108_u0=1'h0;
wire		equals_u90;
wire signed	[31:0]	equals_u90_a_signed;
wire signed	[31:0]	equals_u90_b_signed;
wire		not_u318_u0;
wire		and_u1639_u0;
wire		and_u1640_u0;
wire		and_u1641_u0;
wire		not_u319_u0;
wire		and_u1642_u0;
wire		andOp_u110;
wire		and_u1643_u0;
wire		and_u1644_u0;
wire		not_u320_u0;
wire		simplePinWrite_u287;
wire		or_u444_u0;
reg		reg_0ef045f7_u0=1'h0;
wire		and_u1645_u0;
reg		reg_1ba6eff0_u0=1'h0;
wire		and_u1646_u0;
reg		and_delayed_u109_u0=1'h0;
wire		not_u321_u0;
wire		and_u1647_u0;
wire		and_u1648_u0;
wire		and_u1649_u0;
wire		and_u1650_u0;
wire		not_u322_u0;
wire		simplePinWrite_u288;
wire		and_u1651_u0;
reg		reg_6c316498_u0=1'h0;
reg		reg_6deba007_u0=1'h0;
wire		or_u445_u0;
wire		and_u1652_u0;
reg		reg_2c8794be_u0=1'h0;
reg		and_delayed_u110_u0=1'h0;
wire		and_u1653_u0;
wire		or_u446_u0;
wire		and_u1654_u0;
wire		or_u447_u0;
wire	[1:0]	mux_u156_u0;
reg		and_delayed_u111_u0=1'h0;
wire		and_u1655_u0;
wire		and_u1656_u0;
wire	[1:0]	mux_u157_u0;
wire		or_u448_u0;
wire		or_u449_u0;
wire		or_u450_u0;
wire		and_u1657_u0;
reg		and_delayed_u112_u0=1'h0;
wire		and_u1658_u0;
wire signed	[31:0]	equals_u91_a_signed;
wire		equals_u91;
wire signed	[31:0]	equals_u91_b_signed;
wire		and_u1659_u0;
wire		not_u323_u0;
wire		and_u1660_u0;
wire signed	[31:0]	lessThan_a_signed;
wire		lessThan;
wire signed	[31:0]	lessThan_b_signed;
wire		not_u324_u0;
wire		and_u1661_u0;
wire		and_u1662_u0;
wire		and_u1663_u0;
wire		not_u325_u0;
wire		and_u1664_u0;
wire		simplePinWrite_u289;
wire	[31:0]	add;
reg		reg_62523461_u0=1'h0;
wire		or_u451_u0;
wire		and_u1665_u0;
wire	[31:0]	add_u59;
reg	[15:0]	syncEnable_u153=16'h0;
wire	[15:0]	mux_u158_u0;
reg		reg_4853ac97_u0=1'h0;
wire		and_u1666_u0;
reg	[15:0]	syncEnable_u154_u0=16'h0;
wire		and_u1667_u0;
reg		and_delayed_u113_u0=1'h0;
reg	[2:0]	syncEnable_u155_u0=3'h0;
reg	[15:0]	syncEnable_u156_u0=16'h0;
reg		reg_31498b4c_u0=1'h0;
reg		reg_1f7d581a_u0=1'h0;
wire		and_u1668_u0;
wire		and_u1669_u0;
wire	[31:0]	mux_u159_u0;
reg	[31:0]	syncEnable_u157_u0=32'h0;
wire	[15:0]	mux_u160_u0;
wire		and_u1670_u0;
reg		and_delayed_u114_u0=1'h0;
reg	[31:0]	syncEnable_u158_u0=32'h0;
reg	[15:0]	syncEnable_u159_u0=16'h0;
wire	[31:0]	mux_u161_u0;
wire	[15:0]	mux_u162_u0;
wire		and_u1671_u0;
reg		and_delayed_u115_u0=1'h0;
reg		scoreboard_77421bc3_reg0=1'h0;
reg		scoreboard_77421bc3_reg1=1'h0;
wire		scoreboard_77421bc3_resOr2;
wire		scoreboard_77421bc3_resOr1;
wire		bus_21dc3aa7_;
reg		scoreboard_77421bc3_reg2=1'h0;
wire		scoreboard_77421bc3_and;
wire		scoreboard_77421bc3_resOr0;
wire	[1:0]	mux_u163_u0;
wire		or_u452_u0;
wire		or_u453_u0;
wire	[31:0]	mux_u164_u0;
wire	[31:0]	latch_32d2633c_out;
reg	[31:0]	latch_32d2633c_reg=32'h0;
wire	[31:0]	mux_u165_u0;
wire		or_u454_u0;
reg	[15:0]	latch_19a22e2d_reg=16'h0;
wire	[15:0]	latch_19a22e2d_out;
reg		block_GO_delayed_u4=1'h0;
wire		or_u455_u0;
wire	[1:0]	mux_u166_u0;
reg	[2:0]	syncEnable_u160_u0=3'h0;
reg	[31:0]	syncEnable_u161_u0=32'h0;
reg	[31:0]	syncEnable_u162_u0=32'h0;
reg	[31:0]	syncEnable_u163_u0=32'h0;
reg		block_GO_delayed_u5_u0=1'h0;
reg		syncEnable_u164_u0=1'h0;
reg		syncEnable_u165_u0=1'h0;
reg		syncEnable_u166_u0=1'h0;
reg		syncEnable_u167_u0=1'h0;
reg	[15:0]	syncEnable_u168_u0=16'h0;
reg		syncEnable_u169_u0=1'h0;
reg		syncEnable_u170_u0=1'h0;
wire		and_u1672_u0;
wire	[31:0]	mux_u167_u0;
reg	[15:0]	fbReg_In1Portvalue_u2=16'h0;
reg	[31:0]	fbReg_temp_fsmOldState_LL2_iunzip_2_u0=32'h0;
wire		or_u456_u0;
wire	[15:0]	mux_u168_u0;
reg		loopControl_u2=1'h0;
reg		syncEnable_u171_u0=1'h0;
wire		or_u457_u0;
wire	[31:0]	mux_u169_u0;
reg		reg_68aa9635_u0=1'h0;
wire	[1:0]	mux_u170_u0;
wire		or_u458_u0;
reg		reg_68aa9635_result_delayed_u0=1'h0;
wire		or_u459_u0;
wire	[1:0]	mux_u171_u0;
wire		or_u460_u0;
wire	[31:0]	mux_u172_u0;
wire		mux_u173_u0;
wire		or_u461_u0;
assign equals_a_signed=port_0cb02262_;
assign equals_b_signed=32'h4000;
assign equals=equals_a_signed==equals_b_signed;
assign equals_u86_a_signed=port_0cb02262_;
assign equals_u86_b_signed=32'h4000;
assign equals_u86=equals_u86_a_signed==equals_u86_b_signed;
assign equals_u87_a_signed=port_2710208c_;
assign equals_u87_b_signed=32'h2;
assign equals_u87=equals_u87_a_signed==equals_u87_b_signed;
assign equals_u88_a_signed={30'b0, syncEnable_u160_u0[1:0]};
assign equals_u88_b_signed=32'h0;
assign equals_u88=equals_u88_a_signed==equals_u88_b_signed;
assign not_u311_u0=~equals_u88;
assign and_u1611_u0=block_GO_delayed_u5_u0&equals_u88;
assign and_u1612_u0=block_GO_delayed_u5_u0&not_u311_u0;
assign and_u1613_u0=and_u1618_u0&not_u312_u0;
assign not_u312_u0=~syncEnable_u169_u0;
assign and_u1614_u0=and_u1618_u0&syncEnable_u169_u0;
assign simplePinWrite=and_u1615_u0&{1{and_u1615_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_077142d5_u0<=1'h0;
else reg_077142d5_u0<=reg_2f7b9f51_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_077142d5_result_delayed_u0<=1'h0;
else reg_077142d5_result_delayed_u0<=reg_077142d5_u0;
end
assign or_u434_u0=and_delayed_u103|reg_077142d5_result_delayed_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2f7b9f51_u0<=1'h0;
else reg_2f7b9f51_u0<=and_u1615_u0;
end
assign mux_u153=(and_u1615_u0)?2'h1:2'h3;
assign or_u435_u0=and_u1615_u0|and_u1616_u0;
assign and_u1615_u0=and_u1614_u0&and_u1618_u0;
assign and_u1616_u0=and_u1613_u0&and_u1618_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u103<=1'h0;
else and_delayed_u103<=and_u1616_u0;
end
assign and_u1617_u0=and_u1612_u0&block_GO_delayed_u5_u0;
assign and_u1618_u0=and_u1611_u0&block_GO_delayed_u5_u0;
assign or_u436_u0=or_u434_u0|and_delayed_u104_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u104_u0<=1'h0;
else and_delayed_u104_u0<=and_u1617_u0;
end
assign equals_u89_a_signed={30'b0, syncEnable_u160_u0[1:0]};
assign equals_u89_b_signed=32'h1;
assign equals_u89=equals_u89_a_signed==equals_u89_b_signed;
assign and_u1619_u0=block_GO_delayed_u5_u0&equals_u89;
assign not_u313_u0=~equals_u89;
assign and_u1620_u0=block_GO_delayed_u5_u0&not_u313_u0;
assign and_u1621_u0=and_u1638_u0&syncEnable_u170_u0;
assign and_u1622_u0=and_u1638_u0&not_u314_u0;
assign not_u314_u0=~syncEnable_u170_u0;
assign andOp=port_3777dab3_&port_4cbbb047_;
assign and_u1623_u0=and_u1636_u0&andOp;
assign and_u1624_u0=and_u1636_u0&not_u315_u0;
assign not_u315_u0=~andOp;
assign simplePinWrite_u285=and_u1626_u0&{1{and_u1626_u0}};
assign and_u1625_u0=and_u1624_u0&and_u1636_u0;
assign or_u437_u0=reg_71668bce_u0|and_delayed_u105_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_71668bce_u0<=1'h0;
else reg_71668bce_u0<=reg_76959641_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_76959641_u0<=1'h0;
else reg_76959641_u0<=and_u1626_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u105_u0<=1'h0;
else and_delayed_u105_u0<=and_u1625_u0;
end
assign and_u1626_u0=and_u1623_u0&and_u1636_u0;
assign and_u1627_u0=and_u1635_u0&syncEnable_u164_u0;
assign and_u1628_u0=and_u1635_u0&not_u316_u0;
assign not_u316_u0=~syncEnable_u164_u0;
assign and_u1629_u0=and_u1634_u0&port_4cbbb047_;
assign not_u317_u0=~port_4cbbb047_;
assign and_u1630_u0=and_u1634_u0&not_u317_u0;
assign simplePinWrite_u286=and_u1631_u0&{1{and_u1631_u0}};
assign or_u438_u0=reg_7e4e1b1e_u0|reg_154898a9_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_154898a9_u0<=1'h0;
else reg_154898a9_u0<=and_u1632_u0;
end
assign and_u1631_u0=and_u1629_u0&and_u1634_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u106_u0<=1'h0;
else and_delayed_u106_u0<=and_u1631_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7e4e1b1e_u0<=1'h0;
else reg_7e4e1b1e_u0<=and_delayed_result_delayed_u8;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_result_delayed_u8<=1'h0;
else and_delayed_result_delayed_u8<=and_delayed_u106_u0;
end
assign and_u1632_u0=and_u1630_u0&and_u1634_u0;
assign or_u439_u0=and_u1631_u0|and_u1633_u0;
assign mux_u154_u0=(and_u1631_u0)?2'h2:2'h3;
assign and_u1633_u0=and_u1628_u0&and_u1635_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u107_u0<=1'h0;
else and_delayed_u107_u0<=and_u1633_u0;
end
assign and_u1634_u0=and_u1627_u0&and_u1635_u0;
assign or_u440_u0=or_u438_u0|and_delayed_u107_u0;
assign and_u1635_u0=and_u1622_u0&and_u1638_u0;
assign or_u441_u0=and_u1626_u0|or_u439_u0;
assign mux_u155_u0=(and_u1626_u0)?2'h0:{1'b1, mux_u154_u0[0]};
assign and_u1636_u0=and_u1621_u0&and_u1638_u0;
assign or_u442_u0=or_u437_u0|or_u440_u0;
assign and_u1637_u0=and_u1620_u0&block_GO_delayed_u5_u0;
assign and_u1638_u0=and_u1619_u0&block_GO_delayed_u5_u0;
assign or_u443_u0=or_u442_u0|and_delayed_u108_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u108_u0<=1'h0;
else and_delayed_u108_u0<=and_u1637_u0;
end
assign equals_u90_a_signed={30'b0, syncEnable_u160_u0[1:0]};
assign equals_u90_b_signed=32'h2;
assign equals_u90=equals_u90_a_signed==equals_u90_b_signed;
assign not_u318_u0=~equals_u90;
assign and_u1639_u0=block_GO_delayed_u5_u0&not_u318_u0;
assign and_u1640_u0=block_GO_delayed_u5_u0&equals_u90;
assign and_u1641_u0=and_u1658_u0&syncEnable_u166_u0;
assign not_u319_u0=~syncEnable_u166_u0;
assign and_u1642_u0=and_u1658_u0&not_u319_u0;
assign andOp_u110=port_3777dab3_&port_4cbbb047_;
assign and_u1643_u0=and_u1655_u0&andOp_u110;
assign and_u1644_u0=and_u1655_u0&not_u320_u0;
assign not_u320_u0=~andOp_u110;
assign simplePinWrite_u287=and_u1645_u0&{1{and_u1645_u0}};
assign or_u444_u0=reg_0ef045f7_u0|reg_1ba6eff0_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0ef045f7_u0<=1'h0;
else reg_0ef045f7_u0<=and_delayed_u109_u0;
end
assign and_u1645_u0=and_u1643_u0&and_u1655_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1ba6eff0_u0<=1'h0;
else reg_1ba6eff0_u0<=and_u1646_u0;
end
assign and_u1646_u0=and_u1644_u0&and_u1655_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u109_u0<=1'h0;
else and_delayed_u109_u0<=and_u1645_u0;
end
assign not_u321_u0=~syncEnable_u165_u0;
assign and_u1647_u0=and_u1656_u0&not_u321_u0;
assign and_u1648_u0=and_u1656_u0&syncEnable_u165_u0;
assign and_u1649_u0=and_u1653_u0&not_u322_u0;
assign and_u1650_u0=and_u1653_u0&port_3777dab3_;
assign not_u322_u0=~port_3777dab3_;
assign simplePinWrite_u288=and_u1651_u0&{1{and_u1651_u0}};
assign and_u1651_u0=and_u1650_u0&and_u1653_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6c316498_u0<=1'h0;
else reg_6c316498_u0<=and_u1652_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6deba007_u0<=1'h0;
else reg_6deba007_u0<=reg_2c8794be_u0;
end
assign or_u445_u0=reg_6deba007_u0|reg_6c316498_u0;
assign and_u1652_u0=and_u1649_u0&and_u1653_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2c8794be_u0<=1'h0;
else reg_2c8794be_u0<=and_delayed_u110_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u110_u0<=1'h0;
else and_delayed_u110_u0<=and_u1651_u0;
end
assign and_u1653_u0=and_u1648_u0&and_u1656_u0;
assign or_u446_u0=and_delayed_u111_u0|or_u445_u0;
assign and_u1654_u0=and_u1647_u0&and_u1656_u0;
assign or_u447_u0=and_u1651_u0|and_u1654_u0;
assign mux_u156_u0=(and_u1651_u0)?2'h1:2'h3;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u111_u0<=1'h0;
else and_delayed_u111_u0<=and_u1654_u0;
end
assign and_u1655_u0=and_u1641_u0&and_u1658_u0;
assign and_u1656_u0=and_u1642_u0&and_u1658_u0;
assign mux_u157_u0=(and_u1645_u0)?2'h0:{mux_u156_u0[1], 1'b1};
assign or_u448_u0=and_u1645_u0|or_u447_u0;
assign or_u449_u0=or_u444_u0|or_u446_u0;
assign or_u450_u0=and_delayed_u112_u0|or_u449_u0;
assign and_u1657_u0=and_u1639_u0&block_GO_delayed_u5_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u112_u0<=1'h0;
else and_delayed_u112_u0<=and_u1657_u0;
end
assign and_u1658_u0=and_u1640_u0&block_GO_delayed_u5_u0;
assign equals_u91_a_signed={30'b0, syncEnable_u160_u0[1:0]};
assign equals_u91_b_signed=32'h3;
assign equals_u91=equals_u91_a_signed==equals_u91_b_signed;
assign and_u1659_u0=block_GO_delayed_u5_u0&not_u323_u0;
assign not_u323_u0=~equals_u91;
assign and_u1660_u0=block_GO_delayed_u5_u0&equals_u91;
assign lessThan_a_signed=syncEnable_u161_u0;
assign lessThan_b_signed=syncEnable_u163_u0;
assign lessThan=lessThan_a_signed<lessThan_b_signed;
assign not_u324_u0=~lessThan;
assign and_u1661_u0=and_u1671_u0&not_u324_u0;
assign and_u1662_u0=and_u1671_u0&lessThan;
assign and_u1663_u0=and_u1669_u0&not_u325_u0;
assign not_u325_u0=~syncEnable_u167_u0;
assign and_u1664_u0=and_u1669_u0&syncEnable_u167_u0;
assign simplePinWrite_u289=and_u1667_u0&{1{and_u1667_u0}};
assign add=syncEnable_u161_u0+32'h0;
always @(posedge CLK or posedge and_u1667_u0 or posedge or_u451_u0)
begin
if (or_u451_u0)
reg_62523461_u0<=1'h0;
else if (and_u1667_u0)
reg_62523461_u0<=1'h1;
else reg_62523461_u0<=reg_62523461_u0;
end
assign or_u451_u0=and_u1665_u0|RESET;
assign and_u1665_u0=reg_62523461_u0&port_51623660_;
assign add_u59=syncEnable_u161_u0+32'h1;
always @(posedge CLK)
begin
if (and_u1667_u0)
syncEnable_u153<=port_5a872d3c_;
end
assign mux_u158_u0=(and_delayed_u113_u0)?syncEnable_u154_u0:syncEnable_u153;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4853ac97_u0<=1'h0;
else reg_4853ac97_u0<=and_u1667_u0;
end
assign and_u1666_u0=and_u1663_u0&and_u1669_u0;
always @(posedge CLK)
begin
if (and_u1669_u0)
syncEnable_u154_u0<=syncEnable_u168_u0;
end
assign and_u1667_u0=and_u1664_u0&and_u1669_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u113_u0<=1'h0;
else and_delayed_u113_u0<=and_u1666_u0;
end
always @(posedge CLK)
begin
if (and_u1668_u0)
syncEnable_u155_u0<={1'b0, port_44cbc7ff_};
end
always @(posedge CLK)
begin
if (and_u1671_u0)
syncEnable_u156_u0<=syncEnable_u168_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_31498b4c_u0<=1'h0;
else reg_31498b4c_u0<=and_u1668_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1f7d581a_u0<=1'h0;
else reg_1f7d581a_u0<=and_u1669_u0;
end
assign and_u1668_u0=and_u1661_u0&and_u1671_u0;
assign and_u1669_u0=and_u1662_u0&and_u1671_u0;
assign mux_u159_u0=(reg_1f7d581a_u0)?syncEnable_u157_u0:{30'b0, syncEnable_u155_u0[1:0]};
always @(posedge CLK)
begin
if (and_u1671_u0)
syncEnable_u157_u0<=syncEnable_u162_u0;
end
assign mux_u160_u0=(reg_1f7d581a_u0)?mux_u158_u0:syncEnable_u156_u0;
assign and_u1670_u0=and_u1659_u0&block_GO_delayed_u5_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u114_u0<=1'h0;
else and_delayed_u114_u0<=and_u1670_u0;
end
always @(posedge CLK)
begin
if (block_GO_delayed_u5_u0)
syncEnable_u158_u0<=syncEnable_u162_u0;
end
always @(posedge CLK)
begin
if (block_GO_delayed_u5_u0)
syncEnable_u159_u0<=syncEnable_u168_u0;
end
assign mux_u161_u0=(and_delayed_u115_u0)?mux_u159_u0:syncEnable_u158_u0;
assign mux_u162_u0=(and_delayed_u115_u0)?mux_u160_u0:syncEnable_u159_u0;
assign and_u1671_u0=and_u1660_u0&block_GO_delayed_u5_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u115_u0<=1'h0;
else and_delayed_u115_u0<=and_u1671_u0;
end
always @(posedge CLK)
begin
if (bus_21dc3aa7_)
scoreboard_77421bc3_reg0<=1'h0;
else if (or_u443_u0)
scoreboard_77421bc3_reg0<=1'h1;
else scoreboard_77421bc3_reg0<=scoreboard_77421bc3_reg0;
end
always @(posedge CLK)
begin
if (bus_21dc3aa7_)
scoreboard_77421bc3_reg1<=1'h0;
else if (or_u436_u0)
scoreboard_77421bc3_reg1<=1'h1;
else scoreboard_77421bc3_reg1<=scoreboard_77421bc3_reg1;
end
assign scoreboard_77421bc3_resOr2=or_u450_u0|scoreboard_77421bc3_reg2;
assign scoreboard_77421bc3_resOr1=or_u436_u0|scoreboard_77421bc3_reg1;
assign bus_21dc3aa7_=scoreboard_77421bc3_and|RESET;
always @(posedge CLK)
begin
if (bus_21dc3aa7_)
scoreboard_77421bc3_reg2<=1'h0;
else if (or_u450_u0)
scoreboard_77421bc3_reg2<=1'h1;
else scoreboard_77421bc3_reg2<=scoreboard_77421bc3_reg2;
end
assign scoreboard_77421bc3_and=scoreboard_77421bc3_resOr0&scoreboard_77421bc3_resOr1&scoreboard_77421bc3_resOr2;
assign scoreboard_77421bc3_resOr0=or_u443_u0|scoreboard_77421bc3_reg0;
assign mux_u163_u0=({2{and_u1616_u0}}&2'h0)|({2{and_u1633_u0}}&2'h1)|({2{and_u1654_u0}}&2'h2);
assign or_u452_u0=and_u1616_u0|and_u1633_u0|and_u1654_u0;
assign or_u453_u0=and_u1615_u0|and_u1667_u0;
assign mux_u164_u0=(and_u1615_u0)?32'h0:add_u59;
assign latch_32d2633c_out=(block_GO_delayed_u4)?mux_u161_u0:latch_32d2633c_reg;
always @(posedge CLK)
begin
if (block_GO_delayed_u4)
latch_32d2633c_reg<=mux_u161_u0;
end
assign mux_u165_u0=(and_u1616_u0)?32'h0:32'hfffffffd;
assign or_u454_u0=and_u1616_u0|and_u1668_u0;
always @(posedge CLK)
begin
if (block_GO_delayed_u4)
latch_19a22e2d_reg<=mux_u162_u0;
end
assign latch_19a22e2d_out=(block_GO_delayed_u4)?mux_u162_u0:latch_19a22e2d_reg;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
block_GO_delayed_u4<=1'h0;
else block_GO_delayed_u4<=block_GO_delayed_u5_u0;
end
assign or_u455_u0=or_u435_u0|or_u441_u0|or_u448_u0|and_u1668_u0;
assign mux_u166_u0=({2{or_u435_u0}}&{mux_u153[1], 1'b1})|({2{or_u441_u0}}&mux_u155_u0)|({2{or_u448_u0}}&mux_u157_u0)|({2{and_u1668_u0}}&port_44cbc7ff_);
always @(posedge CLK)
begin
if (and_u1672_u0)
syncEnable_u160_u0<={1'b0, port_57df124f_};
end
always @(posedge CLK)
begin
if (and_u1672_u0)
syncEnable_u161_u0<=port_2710208c_;
end
always @(posedge CLK)
begin
if (and_u1672_u0)
syncEnable_u162_u0<=mux_u167_u0;
end
always @(posedge CLK)
begin
if (and_u1672_u0)
syncEnable_u163_u0<=port_0dedb00e_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
block_GO_delayed_u5_u0<=1'h0;
else block_GO_delayed_u5_u0<=and_u1672_u0;
end
always @(posedge CLK)
begin
if (and_u1672_u0)
syncEnable_u164_u0<=port_2d918d8b_;
end
always @(posedge CLK)
begin
if (and_u1672_u0)
syncEnable_u165_u0<=port_2d918d8b_;
end
always @(posedge CLK)
begin
if (and_u1672_u0)
syncEnable_u166_u0<=equals_u86;
end
always @(posedge CLK)
begin
if (and_u1672_u0)
syncEnable_u167_u0<=port_2d918d8b_;
end
always @(posedge CLK)
begin
if (and_u1672_u0)
syncEnable_u168_u0<=mux_u168_u0;
end
always @(posedge CLK)
begin
if (and_u1672_u0)
syncEnable_u169_u0<=equals_u87;
end
always @(posedge CLK)
begin
if (and_u1672_u0)
syncEnable_u170_u0<=equals;
end
assign and_u1672_u0=or_u456_u0&or_u456_u0;
assign mux_u167_u0=(reg_68aa9635_result_delayed_u0)?32'h0:fbReg_temp_fsmOldState_LL2_iunzip_2_u0;
always @(posedge CLK)
begin
if (scoreboard_77421bc3_and)
fbReg_In1Portvalue_u2<=latch_19a22e2d_out;
end
always @(posedge CLK)
begin
if (scoreboard_77421bc3_and)
fbReg_temp_fsmOldState_LL2_iunzip_2_u0<=latch_32d2633c_out;
end
assign or_u456_u0=reg_68aa9635_result_delayed_u0|loopControl_u2;
assign mux_u168_u0=(reg_68aa9635_result_delayed_u0)?16'h0:fbReg_In1Portvalue_u2;
always @(posedge CLK or posedge syncEnable_u171_u0)
begin
if (syncEnable_u171_u0)
loopControl_u2<=1'h0;
else loopControl_u2<=scoreboard_77421bc3_and;
end
always @(posedge CLK)
begin
if (reg_68aa9635_result_delayed_u0)
syncEnable_u171_u0<=RESET;
end
assign or_u457_u0=GO|or_u454_u0;
assign mux_u169_u0=(GO)?32'hfffffffd:{mux_u165_u0[31:2], 1'b0, mux_u165_u0[0]};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_68aa9635_u0<=1'h0;
else reg_68aa9635_u0<=GO;
end
assign mux_u170_u0=(GO)?2'h0:mux_u163_u0;
assign or_u458_u0=GO|or_u452_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_68aa9635_result_delayed_u0<=1'h0;
else reg_68aa9635_result_delayed_u0<=reg_68aa9635_u0;
end
assign or_u459_u0=GO|or_u455_u0;
assign mux_u171_u0=(GO)?2'h0:mux_u166_u0;
assign or_u460_u0=GO|or_u453_u0;
assign mux_u172_u0=(GO)?32'h0:mux_u164_u0;
assign mux_u173_u0=(GO)?1'h0:1'h1;
assign or_u461_u0=GO|and_u1616_u0;
assign RESULT=or_u458_u0;
assign RESULT_u993=mux_u170_u0;
assign RESULT_u994=or_u459_u0;
assign RESULT_u995=mux_u171_u0;
assign RESULT_u996=or_u460_u0;
assign RESULT_u997=mux_u172_u0;
assign RESULT_u998=or_u457_u0;
assign RESULT_u999={mux_u169_u0[31:2], 1'b0, mux_u169_u0[0]};
assign RESULT_u1000=or_u461_u0;
assign RESULT_u1001=mux_u173_u0;
assign RESULT_u1002=and_u1667_u0;
assign RESULT_u1003=add;
assign RESULT_u1004=port_5a872d3c_;
assign RESULT_u1005=3'h1;
assign RESULT_u1006=simplePinWrite_u287;
assign RESULT_u1007=simplePinWrite_u286;
assign RESULT_u1008=simplePinWrite_u288;
assign RESULT_u1009=simplePinWrite_u289;
assign RESULT_u1010=simplePinWrite;
assign RESULT_u1011=simplePinWrite_u285;
assign DONE=1'h0;
endmodule



module LL2_iunzip_stateVar_In1PortEnable(bus_4b677821_, bus_30c4b424_, bus_2657c6ba_, bus_4371ff51_, bus_6ac01b98_);
input		bus_4b677821_;
input		bus_30c4b424_;
input		bus_2657c6ba_;
input		bus_4371ff51_;
output		bus_6ac01b98_;
reg		stateVar_In1PortEnable_u2=1'h0;
always @(posedge bus_4b677821_ or posedge bus_30c4b424_)
begin
if (bus_30c4b424_)
stateVar_In1PortEnable_u2<=1'h0;
else if (bus_2657c6ba_)
stateVar_In1PortEnable_u2<=bus_4371ff51_;
end
assign bus_6ac01b98_=stateVar_In1PortEnable_u2;
endmodule



module LL2_iunzip_simplememoryreferee_27761197_(bus_60b63314_, bus_0869b5ee_, bus_764c86ba_, bus_43e4e98d_, bus_52c6af95_, bus_524a4e4b_, bus_43a489ea_, bus_5442bd92_, bus_1328384d_, bus_73af1459_, bus_6b014163_, bus_4135f178_, bus_6616c9bf_, bus_188e8a1f_, bus_79e17b19_, bus_055751fe_, bus_5ab9ae07_, bus_3266894e_, bus_4174f34a_, bus_1b8550b0_, bus_7e94d1e2_, bus_0a857fee_, bus_49128048_, bus_098f7792_, bus_1c0ab1f7_, bus_22cdc0fd_, bus_33af47da_, bus_51d68f43_, bus_0e2119bf_);
input		bus_60b63314_;
input		bus_0869b5ee_;
input		bus_764c86ba_;
input	[15:0]	bus_43e4e98d_;
input		bus_52c6af95_;
input	[31:0]	bus_524a4e4b_;
input	[2:0]	bus_43a489ea_;
input		bus_5442bd92_;
input	[31:0]	bus_1328384d_;
input	[2:0]	bus_73af1459_;
input		bus_6b014163_;
input	[31:0]	bus_4135f178_;
input	[2:0]	bus_6616c9bf_;
input		bus_188e8a1f_;
input	[31:0]	bus_79e17b19_;
input	[2:0]	bus_055751fe_;
output	[15:0]	bus_5ab9ae07_;
output	[31:0]	bus_3266894e_;
output		bus_4174f34a_;
output		bus_1b8550b0_;
output	[2:0]	bus_7e94d1e2_;
output	[15:0]	bus_0a857fee_;
output		bus_49128048_;
output	[15:0]	bus_098f7792_;
output		bus_1c0ab1f7_;
output	[15:0]	bus_22cdc0fd_;
output		bus_33af47da_;
output	[15:0]	bus_51d68f43_;
output		bus_0e2119bf_;
wire		not_1bcdba4d_u0;
wire		not_41fe0bfc_u0;
reg		done_qual_u71_u0=1'h0;
wire		and_1c7baefd_u0;
wire		or_0fa8a0a1_u0;
wire		or_5ff43dff_u0;
reg		done_qual_u72_u0=1'h0;
reg		done_qual_u73_u0=1'h0;
wire		not_7bc72bd3_u0;
reg		done_qual_u74_u0=1'h0;
wire		and_060c849a_u0;
wire	[31:0]	mux_374e2914_u0;
wire		or_3168c8f6_u0;
wire		or_7c863926_u0;
wire		and_78a885db_u0;
wire		not_55e397d5_u0;
wire		and_3ef65a8a_u0;
wire		or_40645819_u0;
assign not_1bcdba4d_u0=~bus_764c86ba_;
assign not_41fe0bfc_u0=~bus_764c86ba_;
always @(posedge bus_60b63314_)
begin
if (bus_0869b5ee_)
done_qual_u71_u0<=1'h0;
else done_qual_u71_u0<=bus_188e8a1f_;
end
assign and_1c7baefd_u0=or_5ff43dff_u0&bus_764c86ba_;
assign or_0fa8a0a1_u0=bus_6b014163_|done_qual_u74_u0;
assign or_5ff43dff_u0=bus_5442bd92_|done_qual_u73_u0;
always @(posedge bus_60b63314_)
begin
if (bus_0869b5ee_)
done_qual_u72_u0<=1'h0;
else done_qual_u72_u0<=bus_52c6af95_;
end
always @(posedge bus_60b63314_)
begin
if (bus_0869b5ee_)
done_qual_u73_u0<=1'h0;
else done_qual_u73_u0<=bus_5442bd92_;
end
assign not_7bc72bd3_u0=~bus_764c86ba_;
always @(posedge bus_60b63314_)
begin
if (bus_0869b5ee_)
done_qual_u74_u0<=1'h0;
else done_qual_u74_u0<=bus_6b014163_;
end
assign and_060c849a_u0=or_40645819_u0&bus_764c86ba_;
assign mux_374e2914_u0=({32{bus_52c6af95_}}&bus_524a4e4b_)|({32{bus_5442bd92_}}&bus_1328384d_)|({32{bus_6b014163_}}&bus_4135f178_)|({32{bus_188e8a1f_}}&bus_79e17b19_);
assign or_3168c8f6_u0=bus_52c6af95_|bus_5442bd92_|bus_6b014163_|bus_188e8a1f_;
assign or_7c863926_u0=bus_188e8a1f_|done_qual_u71_u0;
assign bus_5ab9ae07_=16'h0;
assign bus_3266894e_=mux_374e2914_u0;
assign bus_4174f34a_=1'h0;
assign bus_1b8550b0_=or_3168c8f6_u0;
assign bus_7e94d1e2_=3'h1;
assign bus_0a857fee_=bus_43e4e98d_;
assign bus_49128048_=and_060c849a_u0;
assign bus_098f7792_=bus_43e4e98d_;
assign bus_1c0ab1f7_=and_1c7baefd_u0;
assign bus_22cdc0fd_=bus_43e4e98d_;
assign bus_33af47da_=and_3ef65a8a_u0;
assign bus_51d68f43_=bus_43e4e98d_;
assign bus_0e2119bf_=and_78a885db_u0;
assign and_78a885db_u0=or_7c863926_u0&bus_764c86ba_;
assign not_55e397d5_u0=~bus_764c86ba_;
assign and_3ef65a8a_u0=or_0fa8a0a1_u0&bus_764c86ba_;
assign or_40645819_u0=bus_52c6af95_|done_qual_u72_u0;
endmodule



module LL2_iunzip_globalreset_physical_4d3e90cc_(bus_7a7df9cf_, bus_50fc0f9a_, bus_38e1176c_);
input		bus_7a7df9cf_;
input		bus_50fc0f9a_;
output		bus_38e1176c_;
wire		not_4464c834_u0;
reg		glitch_u26=1'h0;
reg		final_u26=1'h1;
wire		or_5c4ce7bb_u0;
reg		cross_u26=1'h0;
reg		sample_u26=1'h0;
wire		and_797ad2e5_u0;
assign not_4464c834_u0=~and_797ad2e5_u0;
always @(posedge bus_7a7df9cf_)
begin
glitch_u26<=cross_u26;
end
always @(posedge bus_7a7df9cf_)
begin
final_u26<=not_4464c834_u0;
end
assign or_5c4ce7bb_u0=bus_50fc0f9a_|final_u26;
assign bus_38e1176c_=or_5c4ce7bb_u0;
always @(posedge bus_7a7df9cf_)
begin
cross_u26<=sample_u26;
end
always @(posedge bus_7a7df9cf_)
begin
sample_u26<=1'h1;
end
assign and_797ad2e5_u0=cross_u26&glitch_u26;
endmodule



module LL2_iunzip_streamFun1(CLK, RESET, GO, port_02b645ca_, port_782b7e63_, port_678d8025_, port_6a7883c4_, port_45c60a90_, port_02d3b259_, port_73617117_, port_32d96ef1_, RESULT, RESULT_u1012, RESULT_u1013, RESULT_u1014, RESULT_u1015, RESULT_u1016, RESULT_u1017, RESULT_u1018, RESULT_u1019, RESULT_u1020, RESULT_u1021, RESULT_u1022, RESULT_u1023, RESULT_u1024, RESULT_u1025, RESULT_u1026, RESULT_u1027, RESULT_u1028, DONE);
input		CLK;
input		RESET;
input		GO;
input		port_02b645ca_;
input	[31:0]	port_782b7e63_;
input		port_678d8025_;
input	[15:0]	port_6a7883c4_;
input		port_45c60a90_;
input	[15:0]	port_02d3b259_;
input		port_73617117_;
input	[15:0]	port_32d96ef1_;
output		RESULT;
output		RESULT_u1012;
output		RESULT_u1013;
output	[31:0]	RESULT_u1014;
output		RESULT_u1015;
output	[31:0]	RESULT_u1016;
output	[2:0]	RESULT_u1017;
output		RESULT_u1018;
output	[31:0]	RESULT_u1019;
output	[2:0]	RESULT_u1020;
output		RESULT_u1021;
output	[31:0]	RESULT_u1022;
output	[15:0]	RESULT_u1023;
output	[2:0]	RESULT_u1024;
output	[15:0]	RESULT_u1025;
output		RESULT_u1026;
output		RESULT_u1027;
output	[15:0]	RESULT_u1028;
output		DONE;
wire		simplePinWrite;
reg		reg_3d761dd7_u0=1'h0;
wire		and_u1674_u0;
wire		or_u462_u0;
wire	[31:0]	add;
wire		and_u1675_u0;
wire	[8:0]	subtract;
wire signed	[8:0]	greaterThanEqualTo_b_signed;
wire		greaterThanEqualTo;
wire signed	[8:0]	greaterThanEqualTo_a_signed;
wire		and_u1676_u0;
wire		not_u326_u0;
wire		and_u1677_u0;
wire	[8:0]	subtract_u16;
wire		and_u1678_u0;
wire		and_u1679_u0;
wire	[8:0]	mux_u174;
wire	[31:0]	add_u60;
wire		and_u1680_u0;
wire		and_u1682_u0;
wire	[16:0]	add_u61;
wire	[15:0]	subtract_u17;
wire	[31:0]	add_u62;
wire		simplePinWrite_u290;
wire	[15:0]	simplePinWrite_u291;
wire	[15:0]	simplePinWrite_u292;
reg	[15:0]	syncEnable_u172=16'h0;
reg	[15:0]	syncEnable_u173_u0=16'h0;
wire	[31:0]	mux_u175_u0;
reg	[15:0]	syncEnable_u174_u0=16'h0;
reg	[31:0]	syncEnable_u175_u0=32'h0;
reg		reg_5f0a2099_u0=1'h0;
reg		reg_0414b780_u0=1'h0;
wire	[31:0]	mux_u176_u0;
wire		or_u463_u0;
reg		reg_5f0a2099_result_delayed_u0=1'h0;
reg	[31:0]	syncEnable_u176_u0=32'h0;
assign simplePinWrite=GO&{1{GO}};
always @(posedge CLK or posedge reg_0414b780_u0 or posedge or_u462_u0)
begin
if (or_u462_u0)
reg_3d761dd7_u0<=1'h0;
else if (reg_0414b780_u0)
reg_3d761dd7_u0<=1'h1;
else reg_3d761dd7_u0<=reg_3d761dd7_u0;
end
assign and_u1674_u0=reg_3d761dd7_u0&port_73617117_;
assign or_u462_u0=and_u1674_u0|RESET;
assign add={31'b0, port_02b645ca_}+32'h0;
assign and_u1675_u0=reg_5f0a2099_u0&port_678d8025_;
assign subtract={8'b0, port_02b645ca_}-9'h1;
assign greaterThanEqualTo_a_signed={subtract[2], subtract[2], subtract[2], subtract[2], subtract[2], subtract[2], subtract[2:0]};
assign greaterThanEqualTo_b_signed=9'h0;
assign greaterThanEqualTo=greaterThanEqualTo_a_signed>=greaterThanEqualTo_b_signed;
assign and_u1676_u0=GO&greaterThanEqualTo;
assign not_u326_u0=~greaterThanEqualTo;
assign and_u1677_u0=GO&not_u326_u0;
assign subtract_u16={8'b0, port_02b645ca_}-9'h1;
assign and_u1678_u0=and_u1676_u0&GO;
assign and_u1679_u0=and_u1677_u0&GO;
assign mux_u174=(and_u1678_u0)?{subtract_u16[2], subtract_u16[2], subtract_u16[2], subtract_u16[2], subtract_u16[2], subtract_u16[2], subtract_u16[2:0]}:9'h2;
assign add_u60={mux_u174[2], mux_u174[2], mux_u174[2], mux_u174[2], mux_u174[2], mux_u174[2], mux_u174[2], mux_u174[2], mux_u174[2], mux_u174[2], mux_u174[2], mux_u174[2], mux_u174[2], mux_u174[2], mux_u174[2], mux_u174[2], mux_u174[2], mux_u174[2], mux_u174[2], mux_u174[2], mux_u174[2], mux_u174[2], mux_u174[2], mux_u174[2], mux_u174[2], mux_u174[2], mux_u174[2], mux_u174[2], mux_u174[2], mux_u174[2:0]}+32'h0;
assign and_u1680_u0=reg_5f0a2099_u0&port_73617117_;
assign and_u1682_u0=reg_5f0a2099_result_delayed_u0&port_678d8025_;
assign add_u61={syncEnable_u174_u0[15], syncEnable_u174_u0}+{port_6a7883c4_[15], port_6a7883c4_};
assign subtract_u17=syncEnable_u172-add_u61[16:1];
assign add_u62=port_782b7e63_+32'h1;
assign simplePinWrite_u290=reg_5f0a2099_result_delayed_u0&{1{reg_5f0a2099_result_delayed_u0}};
assign simplePinWrite_u291=16'h1&{16{1'h1}};
assign simplePinWrite_u292=subtract_u17&{16{reg_5f0a2099_result_delayed_u0}};
always @(posedge CLK)
begin
if (reg_5f0a2099_u0)
syncEnable_u172<=port_6a7883c4_;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u173_u0<=port_32d96ef1_;
end
assign mux_u175_u0=(reg_0414b780_u0)?32'h0:syncEnable_u175_u0;
always @(posedge CLK)
begin
if (reg_5f0a2099_u0)
syncEnable_u174_u0<=port_02d3b259_;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u175_u0<=add_u60;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5f0a2099_u0<=1'h0;
else reg_5f0a2099_u0<=reg_0414b780_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0414b780_u0<=1'h0;
else reg_0414b780_u0<=GO;
end
assign mux_u176_u0=(reg_5f0a2099_u0)?syncEnable_u176_u0:32'h0;
assign or_u463_u0=reg_5f0a2099_u0|reg_5f0a2099_result_delayed_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5f0a2099_result_delayed_u0<=1'h0;
else reg_5f0a2099_result_delayed_u0<=reg_5f0a2099_u0;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u176_u0<={add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2:0]};
end
assign RESULT=GO;
assign RESULT_u1012=1'h0;
assign RESULT_u1013=GO;
assign RESULT_u1014=add_u62;
assign RESULT_u1015=or_u463_u0;
assign RESULT_u1016=mux_u176_u0;
assign RESULT_u1017=3'h1;
assign RESULT_u1018=reg_5f0a2099_u0;
assign RESULT_u1019=mux_u175_u0;
assign RESULT_u1020=3'h1;
assign RESULT_u1021=reg_0414b780_u0;
assign RESULT_u1022=mux_u175_u0;
assign RESULT_u1023=syncEnable_u173_u0;
assign RESULT_u1024=3'h1;
assign RESULT_u1025=simplePinWrite_u292;
assign RESULT_u1026=simplePinWrite_u290;
assign RESULT_u1027=simplePinWrite;
assign RESULT_u1028=simplePinWrite_u291;
assign DONE=reg_5f0a2099_result_delayed_u0;
endmodule



module LL2_iunzip_firstNPixels(CLK, RESET, GO, port_56c10d09_, port_4285ced0_, port_7e889a85_, port_7d5897f1_, port_4bf45ad9_, port_5d69d1a2_, RESULT, RESULT_u1029, RESULT_u1030, RESULT_u1031, RESULT_u1032, RESULT_u1033, RESULT_u1034, RESULT_u1035, RESULT_u1036, RESULT_u1037, RESULT_u1038, RESULT_u1039, DONE);
input		CLK;
input		RESET;
input		GO;
input	[31:0]	port_56c10d09_;
input		port_4285ced0_;
input		port_7e889a85_;
input	[15:0]	port_7d5897f1_;
input		port_4bf45ad9_;
input	[15:0]	port_5d69d1a2_;
output		RESULT;
output	[31:0]	RESULT_u1029;
output		RESULT_u1030;
output	[31:0]	RESULT_u1031;
output	[15:0]	RESULT_u1032;
output	[2:0]	RESULT_u1033;
output		RESULT_u1034;
output	[31:0]	RESULT_u1035;
output	[2:0]	RESULT_u1036;
output		RESULT_u1037;
output	[31:0]	RESULT_u1038;
output	[2:0]	RESULT_u1039;
output		DONE;
wire		and_u1684_u0;
wire		and_u1685_u0;
wire	[31:0]	add;
wire		and_u1686_u0;
wire		or_u464_u0;
reg		reg_03e6937f_u0=1'h0;
wire		or_u465_u0;
reg		reg_1142b8a6_u0=1'h0;
wire		and_u1687_u0;
reg		reg_4025556f_u0=1'h0;
reg	[15:0]	syncEnable_u177=16'h0;
reg		reg_0b5621cb_u0=1'h0;
reg		reg_76aaf2cb_u0=1'h0;
reg	[15:0]	syncEnable_u178_u0=16'h0;
wire		or_u466_u0;
wire	[31:0]	mux_u177;
wire	[15:0]	mux_u178_u0;
assign and_u1684_u0=GO&port_7e889a85_;
assign and_u1685_u0=GO&port_4bf45ad9_;
assign add=port_56c10d09_+32'h2;
assign and_u1686_u0=reg_03e6937f_u0&port_4285ced0_;
assign or_u464_u0=and_u1686_u0|RESET;
always @(posedge CLK or posedge reg_76aaf2cb_u0 or posedge or_u464_u0)
begin
if (or_u464_u0)
reg_03e6937f_u0<=1'h0;
else if (reg_76aaf2cb_u0)
reg_03e6937f_u0<=1'h1;
else reg_03e6937f_u0<=reg_03e6937f_u0;
end
assign or_u465_u0=and_u1687_u0|RESET;
always @(posedge CLK or posedge reg_0b5621cb_u0 or posedge or_u465_u0)
begin
if (or_u465_u0)
reg_1142b8a6_u0<=1'h0;
else if (reg_0b5621cb_u0)
reg_1142b8a6_u0<=1'h1;
else reg_1142b8a6_u0<=reg_1142b8a6_u0;
end
assign and_u1687_u0=reg_1142b8a6_u0&port_4285ced0_;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4025556f_u0<=1'h0;
else reg_4025556f_u0<=reg_0b5621cb_u0;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u177<=port_5d69d1a2_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0b5621cb_u0<=1'h0;
else reg_0b5621cb_u0<=reg_76aaf2cb_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_76aaf2cb_u0<=1'h0;
else reg_76aaf2cb_u0<=GO;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u178_u0<=port_7d5897f1_;
end
assign or_u466_u0=reg_76aaf2cb_u0|reg_0b5621cb_u0;
assign mux_u177=(reg_76aaf2cb_u0)?32'h0:32'h1;
assign mux_u178_u0=(reg_76aaf2cb_u0)?syncEnable_u178_u0:syncEnable_u177;
assign RESULT=GO;
assign RESULT_u1029=add;
assign RESULT_u1030=or_u466_u0;
assign RESULT_u1031={31'b0, mux_u177[0]};
assign RESULT_u1032=mux_u178_u0;
assign RESULT_u1033=3'h1;
assign RESULT_u1034=GO;
assign RESULT_u1035=32'h0;
assign RESULT_u1036=3'h1;
assign RESULT_u1037=GO;
assign RESULT_u1038=32'h1;
assign RESULT_u1039=3'h1;
assign DONE=reg_4025556f_u0;
endmodule



module LL2_iunzip_stateVar_midPoint(bus_68e44dca_, bus_1d3a1112_, bus_0b5520fb_, bus_0cea9df7_, bus_37b6d949_, bus_03a0d5c2_, bus_24329444_, bus_150341ad_, bus_7bdb1d62_, bus_20c3ad1e_, bus_137455cf_);
input		bus_68e44dca_;
input		bus_1d3a1112_;
input		bus_0b5520fb_;
input		bus_0cea9df7_;
input		bus_37b6d949_;
input		bus_03a0d5c2_;
input		bus_24329444_;
input		bus_150341ad_;
input		bus_7bdb1d62_;
input		bus_20c3ad1e_;
output		bus_137455cf_;
reg		stateVar_midPoint_u2=1'h1;
wire		or_12b0b5b9_u0;
always @(posedge bus_68e44dca_ or posedge bus_1d3a1112_)
begin
if (bus_1d3a1112_)
stateVar_midPoint_u2<=1'h1;
else if (or_12b0b5b9_u0)
stateVar_midPoint_u2<=1'h0;
end
assign bus_137455cf_=stateVar_midPoint_u2;
assign or_12b0b5b9_u0=bus_0b5520fb_|bus_37b6d949_|bus_24329444_|bus_7bdb1d62_;
endmodule


