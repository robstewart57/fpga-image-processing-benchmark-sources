// __  ___ __ ___  _ __   ___  ___ 
// \ \/ / '__/ _ \| '_ \ / _ \/ __|
//  >  <| | | (_) | | | | (_) \__ \
// /_/\_\_|  \___/|_| |_|\___/|___/
// 
// Xronos synthesizer version
// Run date: Thu 2 Nov 2017 13:58:38 +0000
// 

module resized_HH1_xy(Out1_COUNT, Out1_RDY, Out1_SEND, Out1_DATA, In1_ACK, In1_COUNT, CLK, RESET, In1_DATA, Out1_ACK, In1_SEND);
output	[15:0]	Out1_COUNT;
input		Out1_RDY;
output		Out1_SEND;
output	[15:0]	Out1_DATA;
output		In1_ACK;
input	[15:0]	In1_COUNT;
wire		reset_go;
wire		repeatRowExpanded_done;
input		CLK;
wire		consumeRow_go;
input		RESET;
wire		reset_done;
input	[15:0]	In1_DATA;
input		Out1_ACK;
wire		repeatRowExpanded_go;
wire		consumeRow_done;
input		In1_SEND;
wire		bus_33b8fb63_;
wire	[15:0]	bus_09fb888a_;
wire		bus_7a2a19b9_;
wire	[15:0]	bus_164dca37_;
wire		bus_7f50b993_;
wire		bus_0b4113f3_;
wire	[15:0]	bus_598e6cc3_;
wire		bus_6e0b18b8_;
wire	[2:0]	bus_639f721f_;
wire	[31:0]	bus_15ad23f9_;
wire	[15:0]	bus_34e7ce30_;
wire		bus_40e60680_;
wire		bus_701b4c75_;
wire		bus_5ddcea96_;
wire		bus_37f5ad72_;
wire	[15:0]	bus_02042397_;
wire	[31:0]	bus_33b10f2a_;
wire		bus_01eb57ef_;
wire	[15:0]	bus_0ed82a61_;
wire	[2:0]	bus_7e23456a_;
wire		bus_6fb584e4_;
wire		bus_393f80fa_;
wire		bus_3a25e3d3_;
wire	[31:0]	bus_45ccd470_;
wire	[31:0]	bus_4159e005_;
wire		bus_02437552_;
wire		resized_HH1_xy_repeatRowExpanded_instance_DONE;
wire	[31:0]	repeatRowExpanded_u5;
wire		repeatRowExpanded_u1;
wire	[31:0]	repeatRowExpanded_u2;
wire	[2:0]	repeatRowExpanded_u7;
wire	[15:0]	repeatRowExpanded_u0;
wire		repeatRowExpanded_u4;
wire	[15:0]	repeatRowExpanded_u6;
wire	[2:0]	repeatRowExpanded_u3;
wire		repeatRowExpanded;
wire		bus_04f762b2_;
wire		resized_HH1_xy_scheduler_instance_DONE;
wire		scheduler_u169;
wire		scheduler_u172;
wire	[31:0]	scheduler_u171;
wire	[15:0]	scheduler_u184;
wire		scheduler_u183;
wire	[15:0]	scheduler_u180;
wire	[31:0]	scheduler_u173;
wire		scheduler_u175;
wire	[31:0]	scheduler_u177;
wire		scheduler_u170;
wire		scheduler_u174;
wire		scheduler_u176;
wire		scheduler_u181;
wire		scheduler;
wire	[31:0]	scheduler_u167;
wire		scheduler_u182;
wire	[2:0]	scheduler_u178;
wire		scheduler_u179;
wire		scheduler_u168;
wire		bus_0ec3b904_;
wire	[15:0]	bus_7b7cec0a_;
wire		resized_HH1_xy_reset_instance_DONE;
wire		reset;
wire	[15:0]	reset_u0;
wire		reset_u1;
wire	[15:0]	reset_u2;
wire		bus_1d017b90_;
wire	[31:0]	bus_7fd1c7f0_;
wire	[15:0]	bus_46857e3b_;
wire	[2:0]	consumeRow_u8;
wire	[2:0]	consumeRow_u4;
wire	[31:0]	consumeRow_u2;
wire		consumeRow_u1;
wire	[15:0]	consumeRow_u3;
wire		consumeRow_u5;
wire		resized_HH1_xy_consumeRow_instance_DONE;
wire	[15:0]	consumeRow_u7;
wire		consumeRow_u9;
wire		consumeRow;
wire	[31:0]	consumeRow_u6;
wire	[15:0]	consumeRow_u0;
wire		bus_652f0115_;
assign Out1_COUNT=scheduler_u180;
assign Out1_SEND=scheduler_u182;
assign Out1_DATA=scheduler_u184;
assign In1_ACK=consumeRow_u9;
assign reset_go=scheduler_u183;
assign repeatRowExpanded_done=bus_652f0115_;
assign consumeRow_go=scheduler_u179;
assign reset_done=bus_0b4113f3_;
assign repeatRowExpanded_go=scheduler_u181;
assign consumeRow_done=bus_7f50b993_;
resized_HH1_xy_Kicker_37 resized_HH1_xy_Kicker_37_1(.CLK(CLK), .RESET(bus_1d017b90_), 
  .bus_33b8fb63_(bus_33b8fb63_));
resized_HH1_xy_structuralmemory_32afea6d_ resized_HH1_xy_structuralmemory_32afea6d__1(.CLK_u8(CLK), 
  .bus_442a9bf6_(bus_1d017b90_), .bus_4a22ea73_(bus_33b10f2a_), .bus_462faa8a_(3'h1), 
  .bus_3de7abb4_(bus_01eb57ef_), .bus_0f5204b8_(bus_37f5ad72_), .bus_30af24a2_(bus_02042397_), 
  .bus_09fb888a_(bus_09fb888a_), .bus_7a2a19b9_(bus_7a2a19b9_));
resized_HH1_xy_stateVar_x resized_HH1_xy_stateVar_x_1(.bus_76da317e_(CLK), .bus_03a06599_(bus_1d017b90_), 
  .bus_356794a6_(consumeRow), .bus_129d31d3_(consumeRow_u0), .bus_34515627_(reset_u1), 
  .bus_5527c111_(16'h0), .bus_164dca37_(bus_164dca37_));
assign bus_7f50b993_=resized_HH1_xy_consumeRow_instance_DONE&{1{resized_HH1_xy_consumeRow_instance_DONE}};
assign bus_0b4113f3_=resized_HH1_xy_reset_instance_DONE&{1{resized_HH1_xy_reset_instance_DONE}};
resized_HH1_xy_simplememoryreferee_69088798_ resized_HH1_xy_simplememoryreferee_69088798__1(.bus_009fa733_(CLK), 
  .bus_735b3be9_(bus_1d017b90_), .bus_100459f6_(bus_0ec3b904_), .bus_74377184_(bus_7b7cec0a_), 
  .bus_4be03c3f_(consumeRow_u1), .bus_26b026db_(consumeRow_u3), .bus_3563aff4_(consumeRow_u2), 
  .bus_7cddbbd4_(3'h1), .bus_4445123e_(repeatRowExpanded_u1), .bus_4d26f206_(repeatRowExpanded_u2), 
  .bus_39458ee1_(3'h1), .bus_598e6cc3_(bus_598e6cc3_), .bus_15ad23f9_(bus_15ad23f9_), 
  .bus_701b4c75_(bus_701b4c75_), .bus_5ddcea96_(bus_5ddcea96_), .bus_639f721f_(bus_639f721f_), 
  .bus_40e60680_(bus_40e60680_), .bus_34e7ce30_(bus_34e7ce30_), .bus_6e0b18b8_(bus_6e0b18b8_));
resized_HH1_xy_simplememoryreferee_7a2b68b8_ resized_HH1_xy_simplememoryreferee_7a2b68b8__1(.bus_3f80456e_(CLK), 
  .bus_4d705476_(bus_1d017b90_), .bus_4c3a3c32_(bus_7a2a19b9_), .bus_35b24d56_(bus_09fb888a_), 
  .bus_02df138a_(consumeRow_u5), .bus_2b98d7b3_(consumeRow_u7), .bus_3cf9cf86_(consumeRow_u6), 
  .bus_2f89026d_(3'h1), .bus_3331e5bc_(repeatRowExpanded_u4), .bus_7ab3b956_(repeatRowExpanded_u6), 
  .bus_72129c42_(repeatRowExpanded_u5), .bus_63363b45_(3'h1), .bus_4ba55bbf_(scheduler_u176), 
  .bus_3bc1a877_(scheduler_u177), .bus_232596ff_(3'h1), .bus_02042397_(bus_02042397_), 
  .bus_33b10f2a_(bus_33b10f2a_), .bus_37f5ad72_(bus_37f5ad72_), .bus_01eb57ef_(bus_01eb57ef_), 
  .bus_7e23456a_(bus_7e23456a_), .bus_6fb584e4_(bus_6fb584e4_), .bus_393f80fa_(bus_393f80fa_), 
  .bus_0ed82a61_(bus_0ed82a61_), .bus_3a25e3d3_(bus_3a25e3d3_));
resized_HH1_xy_stateVar_Out1MaxTokenIndex resized_HH1_xy_stateVar_Out1MaxTokenIndex_1(.bus_5c65caac_(CLK), 
  .bus_70848b9f_(bus_1d017b90_), .bus_602cc7c3_(scheduler_u172), .bus_46e2f861_(scheduler_u173), 
  .bus_45ccd470_(bus_45ccd470_));
resized_HH1_xy_stateVar_fsmOldState_resized_HH1_xy resized_HH1_xy_stateVar_fsmOldState_resized_HH1_xy_1(.bus_1a7328de_(CLK), 
  .bus_33b79498_(bus_1d017b90_), .bus_440ed07c_(scheduler), .bus_48a46ac0_(32'h0), 
  .bus_4159e005_(bus_4159e005_));
resized_HH1_xy_stateVar_Out1PortEnable resized_HH1_xy_stateVar_Out1PortEnable_1(.bus_287bdb2f_(CLK), 
  .bus_65b784d9_(bus_1d017b90_), .bus_461b410b_(scheduler_u174), .bus_690793c8_(scheduler_u175), 
  .bus_02437552_(bus_02437552_));
resized_HH1_xy_repeatRowExpanded resized_HH1_xy_repeatRowExpanded_instance(.CLK(CLK), 
  .RESET(bus_1d017b90_), .GO(repeatRowExpanded_go), .port_0f594897_(bus_46857e3b_), 
  .port_69fc9f4f_(bus_6e0b18b8_), .port_4702c9ee_(bus_34e7ce30_), .port_3b01252b_(bus_393f80fa_), 
  .DONE(resized_HH1_xy_repeatRowExpanded_instance_DONE), .RESULT(repeatRowExpanded), 
  .RESULT_u1075(repeatRowExpanded_u0), .RESULT_u1080(repeatRowExpanded_u1), .RESULT_u1081(repeatRowExpanded_u2), 
  .RESULT_u1082(repeatRowExpanded_u3), .RESULT_u1076(repeatRowExpanded_u4), .RESULT_u1077(repeatRowExpanded_u5), 
  .RESULT_u1078(repeatRowExpanded_u6), .RESULT_u1079(repeatRowExpanded_u7));
resized_HH1_xy_stateVar_fsmState_resized_HH1_xy resized_HH1_xy_stateVar_fsmState_resized_HH1_xy_1(.bus_050f1a62_(CLK), 
  .bus_4af13301_(bus_1d017b90_), .bus_1c39a055_(scheduler_u168), .bus_22b22bb3_(scheduler_u169), 
  .bus_04f762b2_(bus_04f762b2_));
resized_HH1_xy_scheduler resized_HH1_xy_scheduler_instance(.CLK(CLK), .RESET(bus_1d017b90_), 
  .GO(bus_33b8fb63_), .port_57d1c68c_(32'h0), .port_0712fa18_(bus_04f762b2_), .port_5ff18c4c_(bus_7fd1c7f0_), 
  .port_4c4a747e_(bus_45ccd470_), .port_35218c17_(bus_02437552_), .port_0fbd4927_(bus_164dca37_), 
  .port_0d76a61b_(bus_46857e3b_), .port_27356da8_(bus_3a25e3d3_), .port_72850e0c_(bus_0ed82a61_), 
  .port_3599f6c8_(repeatRowExpanded_done), .port_4067da16_(reset_done), .port_6b386c73_(Out1_RDY), 
  .port_67323ff9_(consumeRow_done), .port_316bbc7c_(In1_SEND), .DONE(resized_HH1_xy_scheduler_instance_DONE), 
  .RESULT(scheduler), .RESULT_u1083(scheduler_u167), .RESULT_u1084(scheduler_u168), 
  .RESULT_u1085(scheduler_u169), .RESULT_u1086(scheduler_u170), .RESULT_u1087(scheduler_u171), 
  .RESULT_u1088(scheduler_u172), .RESULT_u1089(scheduler_u173), .RESULT_u1090(scheduler_u174), 
  .RESULT_u1091(scheduler_u175), .RESULT_u1092(scheduler_u176), .RESULT_u1093(scheduler_u177), 
  .RESULT_u1094(scheduler_u178), .RESULT_u1095(scheduler_u179), .RESULT_u1096(scheduler_u180), 
  .RESULT_u1097(scheduler_u181), .RESULT_u1098(scheduler_u182), .RESULT_u1099(scheduler_u183), 
  .RESULT_u1100(scheduler_u184));
resized_HH1_xy_structuralmemory_4abb499d_ resized_HH1_xy_structuralmemory_4abb499d__1(.CLK_u9(CLK), 
  .bus_20b8f358_(bus_1d017b90_), .bus_233a1a3f_(bus_15ad23f9_), .bus_2226f9ce_(3'h1), 
  .bus_7cf55b9c_(bus_5ddcea96_), .bus_5deb4f38_(bus_701b4c75_), .bus_2319feae_(bus_598e6cc3_), 
  .bus_7b7cec0a_(bus_7b7cec0a_), .bus_0ec3b904_(bus_0ec3b904_));
resized_HH1_xy_reset resized_HH1_xy_reset_instance(.CLK(CLK), .RESET(bus_1d017b90_), 
  .GO(reset_go), .DONE(resized_HH1_xy_reset_instance_DONE), .RESULT(reset), .RESULT_u1101(reset_u0), 
  .RESULT_u1102(reset_u1), .RESULT_u1103(reset_u2));
resized_HH1_xy_globalreset_physical_35a1308a_ resized_HH1_xy_globalreset_physical_35a1308a__1(.bus_61966029_(CLK), 
  .bus_12c51121_(RESET), .bus_1d017b90_(bus_1d017b90_));
resized_HH1_xy_stateVar_Out1TokenIndex resized_HH1_xy_stateVar_Out1TokenIndex_1(.bus_4d2a4e2c_(CLK), 
  .bus_65b626e0_(bus_1d017b90_), .bus_4a4819b0_(scheduler_u170), .bus_01d9d88c_(scheduler_u171), 
  .bus_7fd1c7f0_(bus_7fd1c7f0_));
resized_HH1_xy_stateVar_rowRepeated resized_HH1_xy_stateVar_rowRepeated_1(.bus_19552c76_(CLK), 
  .bus_590dd011_(bus_1d017b90_), .bus_52fff2e1_(repeatRowExpanded), .bus_55439b52_(repeatRowExpanded_u0), 
  .bus_6a21e216_(reset), .bus_0bb2ece1_(16'h1), .bus_46857e3b_(bus_46857e3b_));
resized_HH1_xy_consumeRow resized_HH1_xy_consumeRow_instance(.CLK(CLK), .RESET(bus_1d017b90_), 
  .GO(consumeRow_go), .port_531ffb68_(bus_164dca37_), .port_0d7ca19e_(bus_40e60680_), 
  .port_402540c6_(bus_6fb584e4_), .port_2e5e0079_(In1_DATA), .DONE(resized_HH1_xy_consumeRow_instance_DONE), 
  .RESULT(consumeRow), .RESULT_u1104(consumeRow_u0), .RESULT_u1109(consumeRow_u1), 
  .RESULT_u1110(consumeRow_u2), .RESULT_u1111(consumeRow_u3), .RESULT_u1112(consumeRow_u4), 
  .RESULT_u1105(consumeRow_u5), .RESULT_u1106(consumeRow_u6), .RESULT_u1107(consumeRow_u7), 
  .RESULT_u1108(consumeRow_u8), .RESULT_u1113(consumeRow_u9));
assign bus_652f0115_=resized_HH1_xy_repeatRowExpanded_instance_DONE&{1{resized_HH1_xy_repeatRowExpanded_instance_DONE}};
endmodule



module resized_HH1_xy_Kicker_37(CLK, RESET, bus_33b8fb63_);
input		CLK;
input		RESET;
output		bus_33b8fb63_;
reg		kicker_res=1'h0;
wire		bus_597c5469_;
wire		bus_49bdcd82_;
reg		kicker_2=1'h0;
wire		bus_4883aea7_;
reg		kicker_1=1'h0;
wire		bus_3402fa30_;
always @(posedge CLK)
begin
kicker_res<=bus_49bdcd82_;
end
assign bus_597c5469_=bus_3402fa30_&kicker_1;
assign bus_49bdcd82_=kicker_1&bus_3402fa30_&bus_4883aea7_;
always @(posedge CLK)
begin
kicker_2<=bus_597c5469_;
end
assign bus_4883aea7_=~kicker_2;
assign bus_33b8fb63_=kicker_res;
always @(posedge CLK)
begin
kicker_1<=bus_3402fa30_;
end
assign bus_3402fa30_=~RESET;
endmodule



module resized_HH1_xy_forge_memory_512x16_18(CLK, EN, WE, ADDR, DIN, DOUT, DONE);
input		CLK;
input		EN;
input		WE;
input	[31:0]	ADDR;
input	[15:0]	DIN;
output	[15:0]	DOUT;
output		DONE;
wire		we_0;
wire	[15:0]	pre_dout_0;
wire		we_1;
wire	[15:0]	pre_dout_1;
wire		we_2;
wire	[15:0]	pre_dout_2;
wire		we_3;
wire	[15:0]	pre_dout_3;
reg	[15:0]	mux_out;
reg		wen_done;
assign we_0=WE&(ADDR[31:7]==25'h0);
assign we_1=WE&(ADDR[31:7]==25'h1);
assign we_2=WE&(ADDR[31:7]==25'h2);
assign we_3=WE&(ADDR[31:7]==25'h3);
always @(ADDR or pre_dout_0 or pre_dout_1 or pre_dout_2 or pre_dout_3)
begin
case (ADDR[31:7])25'd0:mux_out=pre_dout_0;
25'd1:mux_out=pre_dout_1;
25'd2:mux_out=pre_dout_2;
25'd3:mux_out=pre_dout_3;
default:mux_out=16'h0;
endcase end
always @(posedge CLK)
begin
wen_done<=WE;
end
assign DOUT=mux_out;
assign DONE=EN&!WE|wen_done;
//  Memory array element: COL: 0, ROW: 0
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_0(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[0]), .O(pre_dout_0[0]));
//  Memory array element: COL: 0, ROW: 1
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_1(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[1]), .O(pre_dout_0[1]));
//  Memory array element: COL: 0, ROW: 2
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_2(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[2]), .O(pre_dout_0[2]));
//  Memory array element: COL: 0, ROW: 3
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_3(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[3]), .O(pre_dout_0[3]));
//  Memory array element: COL: 0, ROW: 4
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_4(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[4]), .O(pre_dout_0[4]));
//  Memory array element: COL: 0, ROW: 5
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_5(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[5]), .O(pre_dout_0[5]));
//  Memory array element: COL: 0, ROW: 6
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_6(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[6]), .O(pre_dout_0[6]));
//  Memory array element: COL: 0, ROW: 7
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_7(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[7]), .O(pre_dout_0[7]));
//  Memory array element: COL: 0, ROW: 8
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_8(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[8]), .O(pre_dout_0[8]));
//  Memory array element: COL: 0, ROW: 9
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_9(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[9]), .O(pre_dout_0[9]));
//  Memory array element: COL: 0, ROW: 10
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_10(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[10]), .O(pre_dout_0[10]));
//  Memory array element: COL: 0, ROW: 11
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_11(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[11]), .O(pre_dout_0[11]));
//  Memory array element: COL: 0, ROW: 12
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_12(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[12]), .O(pre_dout_0[12]));
//  Memory array element: COL: 0, ROW: 13
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_13(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[13]), .O(pre_dout_0[13]));
//  Memory array element: COL: 0, ROW: 14
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_14(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[14]), .O(pre_dout_0[14]));
//  Memory array element: COL: 0, ROW: 15
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_15(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[15]), .O(pre_dout_0[15]));
//  Memory array element: COL: 1, ROW: 0
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_16(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[0]), .O(pre_dout_1[0]));
//  Memory array element: COL: 1, ROW: 1
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_17(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[1]), .O(pre_dout_1[1]));
//  Memory array element: COL: 1, ROW: 2
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_18(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[2]), .O(pre_dout_1[2]));
//  Memory array element: COL: 1, ROW: 3
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_19(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[3]), .O(pre_dout_1[3]));
//  Memory array element: COL: 1, ROW: 4
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_20(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[4]), .O(pre_dout_1[4]));
//  Memory array element: COL: 1, ROW: 5
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_21(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[5]), .O(pre_dout_1[5]));
//  Memory array element: COL: 1, ROW: 6
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_22(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[6]), .O(pre_dout_1[6]));
//  Memory array element: COL: 1, ROW: 7
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_23(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[7]), .O(pre_dout_1[7]));
//  Memory array element: COL: 1, ROW: 8
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_24(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[8]), .O(pre_dout_1[8]));
//  Memory array element: COL: 1, ROW: 9
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_25(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[9]), .O(pre_dout_1[9]));
//  Memory array element: COL: 1, ROW: 10
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_26(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[10]), .O(pre_dout_1[10]));
//  Memory array element: COL: 1, ROW: 11
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_27(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[11]), .O(pre_dout_1[11]));
//  Memory array element: COL: 1, ROW: 12
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_28(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[12]), .O(pre_dout_1[12]));
//  Memory array element: COL: 1, ROW: 13
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_29(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[13]), .O(pre_dout_1[13]));
//  Memory array element: COL: 1, ROW: 14
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_30(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[14]), .O(pre_dout_1[14]));
//  Memory array element: COL: 1, ROW: 15
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_31(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[15]), .O(pre_dout_1[15]));
//  Memory array element: COL: 2, ROW: 0
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_32(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[0]), .O(pre_dout_2[0]));
//  Memory array element: COL: 2, ROW: 1
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_33(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[1]), .O(pre_dout_2[1]));
//  Memory array element: COL: 2, ROW: 2
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_34(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[2]), .O(pre_dout_2[2]));
//  Memory array element: COL: 2, ROW: 3
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_35(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[3]), .O(pre_dout_2[3]));
//  Memory array element: COL: 2, ROW: 4
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_36(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[4]), .O(pre_dout_2[4]));
//  Memory array element: COL: 2, ROW: 5
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_37(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[5]), .O(pre_dout_2[5]));
//  Memory array element: COL: 2, ROW: 6
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_38(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[6]), .O(pre_dout_2[6]));
//  Memory array element: COL: 2, ROW: 7
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_39(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[7]), .O(pre_dout_2[7]));
//  Memory array element: COL: 2, ROW: 8
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_40(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[8]), .O(pre_dout_2[8]));
//  Memory array element: COL: 2, ROW: 9
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_41(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[9]), .O(pre_dout_2[9]));
//  Memory array element: COL: 2, ROW: 10
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_42(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[10]), .O(pre_dout_2[10]));
//  Memory array element: COL: 2, ROW: 11
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_43(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[11]), .O(pre_dout_2[11]));
//  Memory array element: COL: 2, ROW: 12
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_44(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[12]), .O(pre_dout_2[12]));
//  Memory array element: COL: 2, ROW: 13
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_45(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[13]), .O(pre_dout_2[13]));
//  Memory array element: COL: 2, ROW: 14
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_46(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[14]), .O(pre_dout_2[14]));
//  Memory array element: COL: 2, ROW: 15
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_47(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[15]), .O(pre_dout_2[15]));
//  Memory array element: COL: 3, ROW: 0
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_48(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[0]), .O(pre_dout_3[0]));
//  Memory array element: COL: 3, ROW: 1
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_49(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[1]), .O(pre_dout_3[1]));
//  Memory array element: COL: 3, ROW: 2
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_50(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[2]), .O(pre_dout_3[2]));
//  Memory array element: COL: 3, ROW: 3
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_51(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[3]), .O(pre_dout_3[3]));
//  Memory array element: COL: 3, ROW: 4
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_52(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[4]), .O(pre_dout_3[4]));
//  Memory array element: COL: 3, ROW: 5
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_53(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[5]), .O(pre_dout_3[5]));
//  Memory array element: COL: 3, ROW: 6
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_54(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[6]), .O(pre_dout_3[6]));
//  Memory array element: COL: 3, ROW: 7
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_55(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[7]), .O(pre_dout_3[7]));
//  Memory array element: COL: 3, ROW: 8
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_56(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[8]), .O(pre_dout_3[8]));
//  Memory array element: COL: 3, ROW: 9
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_57(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[9]), .O(pre_dout_3[9]));
//  Memory array element: COL: 3, ROW: 10
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_58(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[10]), .O(pre_dout_3[10]));
//  Memory array element: COL: 3, ROW: 11
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_59(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[11]), .O(pre_dout_3[11]));
//  Memory array element: COL: 3, ROW: 12
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_60(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[12]), .O(pre_dout_3[12]));
//  Memory array element: COL: 3, ROW: 13
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_61(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[13]), .O(pre_dout_3[13]));
//  Memory array element: COL: 3, ROW: 14
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_62(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[14]), .O(pre_dout_3[14]));
//  Memory array element: COL: 3, ROW: 15
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_63(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[15]), .O(pre_dout_3[15]));
endmodule



module resized_HH1_xy_structuralmemory_32afea6d_(CLK_u8, bus_442a9bf6_, bus_4a22ea73_, bus_462faa8a_, bus_3de7abb4_, bus_0f5204b8_, bus_30af24a2_, bus_09fb888a_, bus_7a2a19b9_);
input		CLK_u8;
input		bus_442a9bf6_;
input	[31:0]	bus_4a22ea73_;
input	[2:0]	bus_462faa8a_;
input		bus_3de7abb4_;
input		bus_0f5204b8_;
input	[15:0]	bus_30af24a2_;
output	[15:0]	bus_09fb888a_;
output		bus_7a2a19b9_;
wire		not_764a55cf_u0;
wire	[15:0]	bus_6b50a464_;
reg		logicalMem_4027b80d_we_delay0_u0=1'h0;
wire		or_3b5c7fc0_u0;
wire		or_13d423a9_u0;
wire		and_475306ed_u0;
assign not_764a55cf_u0=~bus_0f5204b8_;
assign bus_09fb888a_=bus_6b50a464_;
assign bus_7a2a19b9_=or_3b5c7fc0_u0;
resized_HH1_xy_forge_memory_512x16_18 resized_HH1_xy_forge_memory_512x16_18_instance0(.CLK(CLK_u8), 
  .EN(or_13d423a9_u0), .WE(bus_0f5204b8_), .ADDR(bus_4a22ea73_), .DIN(bus_30af24a2_), 
  .DOUT(bus_6b50a464_), .DONE());
always @(posedge CLK_u8 or posedge bus_442a9bf6_)
begin
if (bus_442a9bf6_)
logicalMem_4027b80d_we_delay0_u0<=1'h0;
else logicalMem_4027b80d_we_delay0_u0<=bus_0f5204b8_;
end
assign or_3b5c7fc0_u0=and_475306ed_u0|logicalMem_4027b80d_we_delay0_u0;
assign or_13d423a9_u0=bus_3de7abb4_|bus_0f5204b8_;
assign and_475306ed_u0=bus_3de7abb4_&not_764a55cf_u0;
endmodule



module resized_HH1_xy_endianswapper_7b71ad0a_(endianswapper_7b71ad0a_in, endianswapper_7b71ad0a_out);
input	[15:0]	endianswapper_7b71ad0a_in;
output	[15:0]	endianswapper_7b71ad0a_out;
assign endianswapper_7b71ad0a_out=endianswapper_7b71ad0a_in;
endmodule



module resized_HH1_xy_endianswapper_18e73629_(endianswapper_18e73629_in, endianswapper_18e73629_out);
input	[15:0]	endianswapper_18e73629_in;
output	[15:0]	endianswapper_18e73629_out;
assign endianswapper_18e73629_out=endianswapper_18e73629_in;
endmodule



module resized_HH1_xy_stateVar_x(bus_76da317e_, bus_03a06599_, bus_356794a6_, bus_129d31d3_, bus_34515627_, bus_5527c111_, bus_164dca37_);
input		bus_76da317e_;
input		bus_03a06599_;
input		bus_356794a6_;
input	[15:0]	bus_129d31d3_;
input		bus_34515627_;
input	[15:0]	bus_5527c111_;
output	[15:0]	bus_164dca37_;
wire	[15:0]	mux_04bad6f0_u0;
wire	[15:0]	endianswapper_7b71ad0a_out;
wire		or_1c2cc8d1_u0;
wire	[15:0]	endianswapper_18e73629_out;
reg	[15:0]	stateVar_x_u0=16'h0;
assign bus_164dca37_=endianswapper_7b71ad0a_out;
assign mux_04bad6f0_u0=(bus_356794a6_)?bus_129d31d3_:16'h0;
resized_HH1_xy_endianswapper_7b71ad0a_ resized_HH1_xy_endianswapper_7b71ad0a__1(.endianswapper_7b71ad0a_in(stateVar_x_u0), 
  .endianswapper_7b71ad0a_out(endianswapper_7b71ad0a_out));
assign or_1c2cc8d1_u0=bus_356794a6_|bus_34515627_;
resized_HH1_xy_endianswapper_18e73629_ resized_HH1_xy_endianswapper_18e73629__1(.endianswapper_18e73629_in(mux_04bad6f0_u0), 
  .endianswapper_18e73629_out(endianswapper_18e73629_out));
always @(posedge bus_76da317e_ or posedge bus_03a06599_)
begin
if (bus_03a06599_)
stateVar_x_u0<=16'h0;
else if (or_1c2cc8d1_u0)
stateVar_x_u0<=endianswapper_18e73629_out;
end
endmodule



module resized_HH1_xy_simplememoryreferee_69088798_(bus_009fa733_, bus_735b3be9_, bus_100459f6_, bus_74377184_, bus_4be03c3f_, bus_26b026db_, bus_3563aff4_, bus_7cddbbd4_, bus_4445123e_, bus_4d26f206_, bus_39458ee1_, bus_598e6cc3_, bus_15ad23f9_, bus_701b4c75_, bus_5ddcea96_, bus_639f721f_, bus_40e60680_, bus_34e7ce30_, bus_6e0b18b8_);
input		bus_009fa733_;
input		bus_735b3be9_;
input		bus_100459f6_;
input	[15:0]	bus_74377184_;
input		bus_4be03c3f_;
input	[15:0]	bus_26b026db_;
input	[31:0]	bus_3563aff4_;
input	[2:0]	bus_7cddbbd4_;
input		bus_4445123e_;
input	[31:0]	bus_4d26f206_;
input	[2:0]	bus_39458ee1_;
output	[15:0]	bus_598e6cc3_;
output	[31:0]	bus_15ad23f9_;
output		bus_701b4c75_;
output		bus_5ddcea96_;
output	[2:0]	bus_639f721f_;
output		bus_40e60680_;
output	[15:0]	bus_34e7ce30_;
output		bus_6e0b18b8_;
wire		and_5745a805_u0;
reg		done_qual_u75=1'h0;
wire	[31:0]	mux_1c38951c_u0;
wire		and_50105215_u0;
wire	[15:0]	mux_0275843a_u0;
reg		done_qual_u76_u0=1'h0;
wire		or_5fc0b6b2_u0;
wire		not_74826954_u0;
wire		or_6ba811b1_u0;
wire		not_323d9867_u0;
wire		or_41b4d4e8_u0;
assign and_5745a805_u0=or_6ba811b1_u0&bus_100459f6_;
always @(posedge bus_009fa733_)
begin
if (bus_735b3be9_)
done_qual_u75<=1'h0;
else done_qual_u75<=bus_4445123e_;
end
assign mux_1c38951c_u0=(bus_4be03c3f_)?bus_3563aff4_:bus_4d26f206_;
assign and_50105215_u0=or_41b4d4e8_u0&bus_100459f6_;
assign mux_0275843a_u0=({16{bus_4be03c3f_}}&bus_26b026db_);
always @(posedge bus_009fa733_)
begin
if (bus_735b3be9_)
done_qual_u76_u0<=1'h0;
else done_qual_u76_u0<=bus_4be03c3f_;
end
assign or_5fc0b6b2_u0=bus_4be03c3f_|bus_4445123e_;
assign not_74826954_u0=~bus_100459f6_;
assign bus_598e6cc3_=mux_0275843a_u0;
assign bus_15ad23f9_=mux_1c38951c_u0;
assign bus_701b4c75_=bus_4be03c3f_;
assign bus_5ddcea96_=or_5fc0b6b2_u0;
assign bus_639f721f_=3'h1;
assign bus_40e60680_=and_50105215_u0;
assign bus_34e7ce30_=bus_74377184_;
assign bus_6e0b18b8_=and_5745a805_u0;
assign or_6ba811b1_u0=bus_4445123e_|done_qual_u75;
assign not_323d9867_u0=~bus_100459f6_;
assign or_41b4d4e8_u0=bus_4be03c3f_|done_qual_u76_u0;
endmodule



module resized_HH1_xy_simplememoryreferee_7a2b68b8_(bus_3f80456e_, bus_4d705476_, bus_4c3a3c32_, bus_35b24d56_, bus_02df138a_, bus_2b98d7b3_, bus_3cf9cf86_, bus_2f89026d_, bus_3331e5bc_, bus_7ab3b956_, bus_72129c42_, bus_63363b45_, bus_4ba55bbf_, bus_3bc1a877_, bus_232596ff_, bus_02042397_, bus_33b10f2a_, bus_37f5ad72_, bus_01eb57ef_, bus_7e23456a_, bus_6fb584e4_, bus_393f80fa_, bus_0ed82a61_, bus_3a25e3d3_);
input		bus_3f80456e_;
input		bus_4d705476_;
input		bus_4c3a3c32_;
input	[15:0]	bus_35b24d56_;
input		bus_02df138a_;
input	[15:0]	bus_2b98d7b3_;
input	[31:0]	bus_3cf9cf86_;
input	[2:0]	bus_2f89026d_;
input		bus_3331e5bc_;
input	[15:0]	bus_7ab3b956_;
input	[31:0]	bus_72129c42_;
input	[2:0]	bus_63363b45_;
input		bus_4ba55bbf_;
input	[31:0]	bus_3bc1a877_;
input	[2:0]	bus_232596ff_;
output	[15:0]	bus_02042397_;
output	[31:0]	bus_33b10f2a_;
output		bus_37f5ad72_;
output		bus_01eb57ef_;
output	[2:0]	bus_7e23456a_;
output		bus_6fb584e4_;
output		bus_393f80fa_;
output	[15:0]	bus_0ed82a61_;
output		bus_3a25e3d3_;
wire		not_5a672cc6_u0;
reg		done_qual_u77_u0=1'h0;
wire		or_4a25d061_u0;
wire		or_449bd1dc_u0;
wire		or_249c3116_u0;
wire		or_6d1c2ccc_u0;
wire		or_32ea375b_u0;
wire		not_29b40485_u0;
wire		not_23801f91_u0;
wire	[15:0]	mux_50fa2648_u0;
wire		and_0b9ae0a9_u0;
reg		done_qual_u78_u0=1'h0;
wire		and_4207ed7e_u0;
wire		and_04ef60b1_u0;
wire	[31:0]	mux_1d2a54b5_u0;
reg		done_qual_u79_u0=1'h0;
assign not_5a672cc6_u0=~bus_4c3a3c32_;
always @(posedge bus_3f80456e_)
begin
if (bus_4d705476_)
done_qual_u77_u0<=1'h0;
else done_qual_u77_u0<=bus_4ba55bbf_;
end
assign or_4a25d061_u0=bus_4ba55bbf_|done_qual_u77_u0;
assign or_449bd1dc_u0=bus_02df138a_|bus_3331e5bc_;
assign bus_02042397_=mux_50fa2648_u0;
assign bus_33b10f2a_=mux_1d2a54b5_u0;
assign bus_37f5ad72_=or_449bd1dc_u0;
assign bus_01eb57ef_=or_6d1c2ccc_u0;
assign bus_7e23456a_=3'h1;
assign bus_6fb584e4_=and_4207ed7e_u0;
assign bus_393f80fa_=and_04ef60b1_u0;
assign bus_0ed82a61_=bus_35b24d56_;
assign bus_3a25e3d3_=and_0b9ae0a9_u0;
assign or_249c3116_u0=bus_3331e5bc_|done_qual_u79_u0;
assign or_6d1c2ccc_u0=bus_02df138a_|bus_3331e5bc_|bus_4ba55bbf_;
assign or_32ea375b_u0=bus_02df138a_|done_qual_u78_u0;
assign not_29b40485_u0=~bus_4c3a3c32_;
assign not_23801f91_u0=~bus_4c3a3c32_;
assign mux_50fa2648_u0=(bus_02df138a_)?bus_2b98d7b3_:bus_7ab3b956_;
assign and_0b9ae0a9_u0=or_4a25d061_u0&bus_4c3a3c32_;
always @(posedge bus_3f80456e_)
begin
if (bus_4d705476_)
done_qual_u78_u0<=1'h0;
else done_qual_u78_u0<=bus_02df138a_;
end
assign and_4207ed7e_u0=or_32ea375b_u0&bus_4c3a3c32_;
assign and_04ef60b1_u0=or_249c3116_u0&bus_4c3a3c32_;
assign mux_1d2a54b5_u0=({32{bus_02df138a_}}&bus_3cf9cf86_)|({32{bus_3331e5bc_}}&bus_72129c42_)|({32{bus_4ba55bbf_}}&bus_3bc1a877_);
always @(posedge bus_3f80456e_)
begin
if (bus_4d705476_)
done_qual_u79_u0<=1'h0;
else done_qual_u79_u0<=bus_3331e5bc_;
end
endmodule



module resized_HH1_xy_endianswapper_0096a48d_(endianswapper_0096a48d_in, endianswapper_0096a48d_out);
input	[31:0]	endianswapper_0096a48d_in;
output	[31:0]	endianswapper_0096a48d_out;
assign endianswapper_0096a48d_out=endianswapper_0096a48d_in;
endmodule



module resized_HH1_xy_endianswapper_086443cf_(endianswapper_086443cf_in, endianswapper_086443cf_out);
input	[31:0]	endianswapper_086443cf_in;
output	[31:0]	endianswapper_086443cf_out;
assign endianswapper_086443cf_out=endianswapper_086443cf_in;
endmodule



module resized_HH1_xy_stateVar_Out1MaxTokenIndex(bus_5c65caac_, bus_70848b9f_, bus_602cc7c3_, bus_46e2f861_, bus_45ccd470_);
input		bus_5c65caac_;
input		bus_70848b9f_;
input		bus_602cc7c3_;
input	[31:0]	bus_46e2f861_;
output	[31:0]	bus_45ccd470_;
wire	[31:0]	endianswapper_0096a48d_out;
wire	[31:0]	endianswapper_086443cf_out;
reg	[31:0]	stateVar_Out1MaxTokenIndex_u0=32'h0;
assign bus_45ccd470_=endianswapper_086443cf_out;
resized_HH1_xy_endianswapper_0096a48d_ resized_HH1_xy_endianswapper_0096a48d__1(.endianswapper_0096a48d_in(bus_46e2f861_), 
  .endianswapper_0096a48d_out(endianswapper_0096a48d_out));
resized_HH1_xy_endianswapper_086443cf_ resized_HH1_xy_endianswapper_086443cf__1(.endianswapper_086443cf_in(stateVar_Out1MaxTokenIndex_u0), 
  .endianswapper_086443cf_out(endianswapper_086443cf_out));
always @(posedge bus_5c65caac_ or posedge bus_70848b9f_)
begin
if (bus_70848b9f_)
stateVar_Out1MaxTokenIndex_u0<=32'h0;
else if (bus_602cc7c3_)
stateVar_Out1MaxTokenIndex_u0<=endianswapper_0096a48d_out;
end
endmodule



module resized_HH1_xy_endianswapper_462ffbdd_(endianswapper_462ffbdd_in, endianswapper_462ffbdd_out);
input	[31:0]	endianswapper_462ffbdd_in;
output	[31:0]	endianswapper_462ffbdd_out;
assign endianswapper_462ffbdd_out=32'h0;
endmodule



module resized_HH1_xy_endianswapper_6e5c7ccb_(endianswapper_6e5c7ccb_in, endianswapper_6e5c7ccb_out);
input	[31:0]	endianswapper_6e5c7ccb_in;
output	[31:0]	endianswapper_6e5c7ccb_out;
assign endianswapper_6e5c7ccb_out=32'h0;
endmodule



module resized_HH1_xy_stateVar_fsmOldState_resized_HH1_xy(bus_1a7328de_, bus_33b79498_, bus_440ed07c_, bus_48a46ac0_, bus_4159e005_);
input		bus_1a7328de_;
input		bus_33b79498_;
input		bus_440ed07c_;
input	[31:0]	bus_48a46ac0_;
output	[31:0]	bus_4159e005_;
wire	[31:0]	endianswapper_462ffbdd_out;
wire	[31:0]	endianswapper_6e5c7ccb_out;
resized_HH1_xy_endianswapper_462ffbdd_ resized_HH1_xy_endianswapper_462ffbdd__1(.endianswapper_462ffbdd_in(32'h0), 
  .endianswapper_462ffbdd_out(endianswapper_462ffbdd_out));
assign bus_4159e005_=32'h0;
resized_HH1_xy_endianswapper_6e5c7ccb_ resized_HH1_xy_endianswapper_6e5c7ccb__1(.endianswapper_6e5c7ccb_in(32'h0), 
  .endianswapper_6e5c7ccb_out(endianswapper_6e5c7ccb_out));
endmodule



module resized_HH1_xy_stateVar_Out1PortEnable(bus_287bdb2f_, bus_65b784d9_, bus_461b410b_, bus_690793c8_, bus_02437552_);
input		bus_287bdb2f_;
input		bus_65b784d9_;
input		bus_461b410b_;
input		bus_690793c8_;
output		bus_02437552_;
reg		stateVar_Out1PortEnable_u0=1'h0;
assign bus_02437552_=stateVar_Out1PortEnable_u0;
always @(posedge bus_287bdb2f_ or posedge bus_65b784d9_)
begin
if (bus_65b784d9_)
stateVar_Out1PortEnable_u0<=1'h0;
else if (bus_461b410b_)
stateVar_Out1PortEnable_u0<=bus_690793c8_;
end
endmodule



module resized_HH1_xy_repeatRowExpanded(CLK, RESET, GO, port_0f594897_, port_3b01252b_, port_69fc9f4f_, port_4702c9ee_, RESULT, RESULT_u1075, RESULT_u1076, RESULT_u1077, RESULT_u1078, RESULT_u1079, RESULT_u1080, RESULT_u1081, RESULT_u1082, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_0f594897_;
input		port_3b01252b_;
input		port_69fc9f4f_;
input	[15:0]	port_4702c9ee_;
output		RESULT;
output	[15:0]	RESULT_u1075;
output		RESULT_u1076;
output	[31:0]	RESULT_u1077;
output	[15:0]	RESULT_u1078;
output	[2:0]	RESULT_u1079;
output		RESULT_u1080;
output	[31:0]	RESULT_u1081;
output	[2:0]	RESULT_u1082;
output		DONE;
wire	[15:0]	add;
wire	[31:0]	add_u65;
wire		and_u1748_u0;
wire	[31:0]	add_u66;
wire		and_u1749_u0;
wire		or_u479_u0;
reg		reg_6b6ad240_u0=1'h0;
wire	[31:0]	add_u67;
reg	[31:0]	syncEnable_u179=32'h0;
wire signed	[31:0]	lessThan_b_signed;
wire		lessThan;
wire signed	[31:0]	lessThan_a_signed;
wire		and_u1750_u0;
wire		not_u345_u0;
wire		and_u1751_u0;
reg		reg_75530b9a_u0=1'h0;
wire		and_u1752_u0;
wire		and_u1753_u0;
wire	[31:0]	mux_u179;
wire		or_u480_u0;
reg		reg_6d2a7e38_u0=1'h0;
assign add=port_0f594897_+16'h1;
assign add_u65=mux_u179+32'h0;
assign and_u1748_u0=and_u1752_u0&port_69fc9f4f_;
assign add_u66=mux_u179+32'h0;
assign and_u1749_u0=reg_6b6ad240_u0&port_3b01252b_;
assign or_u479_u0=and_u1749_u0|RESET;
always @(posedge CLK or posedge and_u1752_u0 or posedge or_u479_u0)
begin
if (or_u479_u0)
reg_6b6ad240_u0<=1'h0;
else if (and_u1752_u0)
reg_6b6ad240_u0<=1'h1;
else reg_6b6ad240_u0<=reg_6b6ad240_u0;
end
assign add_u67=mux_u179+32'h1;
always @(posedge CLK)
begin
if (and_u1752_u0)
syncEnable_u179<=add_u67;
end
assign lessThan_a_signed=mux_u179;
assign lessThan_b_signed=32'h200;
assign lessThan=lessThan_a_signed<lessThan_b_signed;
assign and_u1750_u0=or_u480_u0&not_u345_u0;
assign not_u345_u0=~lessThan;
assign and_u1751_u0=or_u480_u0&lessThan;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_75530b9a_u0<=1'h0;
else reg_75530b9a_u0<=and_u1752_u0;
end
assign and_u1752_u0=and_u1751_u0&or_u480_u0;
assign and_u1753_u0=and_u1750_u0&or_u480_u0;
assign mux_u179=(reg_6d2a7e38_u0)?32'h0:syncEnable_u179;
assign or_u480_u0=reg_6d2a7e38_u0|reg_75530b9a_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6d2a7e38_u0<=1'h0;
else reg_6d2a7e38_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u1075=add;
assign RESULT_u1076=and_u1752_u0;
assign RESULT_u1077=add_u66;
assign RESULT_u1078=port_4702c9ee_;
assign RESULT_u1079=3'h1;
assign RESULT_u1080=and_u1752_u0;
assign RESULT_u1081=add_u65;
assign RESULT_u1082=3'h1;
assign DONE=and_u1753_u0;
endmodule



module resized_HH1_xy_endianswapper_17cc46ad_(endianswapper_17cc46ad_in, endianswapper_17cc46ad_out);
input		endianswapper_17cc46ad_in;
output		endianswapper_17cc46ad_out;
assign endianswapper_17cc46ad_out=endianswapper_17cc46ad_in;
endmodule



module resized_HH1_xy_endianswapper_688d46be_(endianswapper_688d46be_in, endianswapper_688d46be_out);
input		endianswapper_688d46be_in;
output		endianswapper_688d46be_out;
assign endianswapper_688d46be_out=endianswapper_688d46be_in;
endmodule



module resized_HH1_xy_stateVar_fsmState_resized_HH1_xy(bus_050f1a62_, bus_4af13301_, bus_1c39a055_, bus_22b22bb3_, bus_04f762b2_);
input		bus_050f1a62_;
input		bus_4af13301_;
input		bus_1c39a055_;
input		bus_22b22bb3_;
output		bus_04f762b2_;
wire		endianswapper_17cc46ad_out;
wire		endianswapper_688d46be_out;
reg		stateVar_fsmState_resized_HH1_xy_u0=1'h0;
resized_HH1_xy_endianswapper_17cc46ad_ resized_HH1_xy_endianswapper_17cc46ad__1(.endianswapper_17cc46ad_in(stateVar_fsmState_resized_HH1_xy_u0), 
  .endianswapper_17cc46ad_out(endianswapper_17cc46ad_out));
resized_HH1_xy_endianswapper_688d46be_ resized_HH1_xy_endianswapper_688d46be__1(.endianswapper_688d46be_in(bus_22b22bb3_), 
  .endianswapper_688d46be_out(endianswapper_688d46be_out));
always @(posedge bus_050f1a62_ or posedge bus_4af13301_)
begin
if (bus_4af13301_)
stateVar_fsmState_resized_HH1_xy_u0<=1'h0;
else if (bus_1c39a055_)
stateVar_fsmState_resized_HH1_xy_u0<=endianswapper_688d46be_out;
end
assign bus_04f762b2_=endianswapper_17cc46ad_out;
endmodule



module resized_HH1_xy_scheduler(CLK, RESET, GO, port_57d1c68c_, port_0712fa18_, port_5ff18c4c_, port_4c4a747e_, port_35218c17_, port_0fbd4927_, port_0d76a61b_, port_27356da8_, port_72850e0c_, port_3599f6c8_, port_4067da16_, port_6b386c73_, port_67323ff9_, port_316bbc7c_, RESULT, RESULT_u1083, RESULT_u1084, RESULT_u1085, RESULT_u1086, RESULT_u1087, RESULT_u1088, RESULT_u1089, RESULT_u1090, RESULT_u1091, RESULT_u1092, RESULT_u1093, RESULT_u1094, RESULT_u1095, RESULT_u1096, RESULT_u1097, RESULT_u1098, RESULT_u1099, RESULT_u1100, DONE);
input		CLK;
input		RESET;
input		GO;
input	[31:0]	port_57d1c68c_;
input		port_0712fa18_;
input	[31:0]	port_5ff18c4c_;
input	[31:0]	port_4c4a747e_;
input		port_35218c17_;
input	[15:0]	port_0fbd4927_;
input	[15:0]	port_0d76a61b_;
input		port_27356da8_;
input	[15:0]	port_72850e0c_;
input		port_3599f6c8_;
input		port_4067da16_;
input		port_6b386c73_;
input		port_67323ff9_;
input		port_316bbc7c_;
output		RESULT;
output	[31:0]	RESULT_u1083;
output		RESULT_u1084;
output		RESULT_u1085;
output		RESULT_u1086;
output	[31:0]	RESULT_u1087;
output		RESULT_u1088;
output	[31:0]	RESULT_u1089;
output		RESULT_u1090;
output		RESULT_u1091;
output		RESULT_u1092;
output	[31:0]	RESULT_u1093;
output	[2:0]	RESULT_u1094;
output		RESULT_u1095;
output	[15:0]	RESULT_u1096;
output		RESULT_u1097;
output		RESULT_u1098;
output		RESULT_u1099;
output	[15:0]	RESULT_u1100;
output		DONE;
wire		and_u1754_u0;
wire	[15:0]	lessThan_a_unsigned;
wire	[15:0]	lessThan_b_unsigned;
wire		lessThan;
wire	[15:0]	equals_a_unsigned;
wire	[15:0]	equals_b_unsigned;
wire		equals;
wire		lessThan_u38;
wire	[15:0]	lessThan_u38_b_unsigned;
wire	[15:0]	lessThan_u38_a_unsigned;
wire		andOp;
wire		equals_u92;
wire	[15:0]	equals_u92_a_unsigned;
wire	[15:0]	equals_u92_b_unsigned;
wire		equals_u93;
wire signed	[31:0]	equals_u93_a_signed;
wire signed	[31:0]	equals_u93_b_signed;
wire		not_u346_u0;
wire		and_u1755_u0;
wire		and_u1756_u0;
wire		andOp_u113;
wire		not_u347_u0;
wire		and_u1757_u0;
wire		and_u1758_u0;
wire		simplePinWrite;
wire		and_u1759_u0;
wire		and_u1760_u0;
wire		not_u348_u0;
wire		simplePinWrite_u316;
wire		and_u1761_u0;
wire		not_u349_u0;
wire		and_u1762_u0;
wire		simplePinWrite_u317;
wire		and_u1763_u0;
reg		reg_608e408d_u0=1'h0;
reg		reg_3d110516_u0=1'h0;
reg		reg_745e0c57_u0=1'h0;
reg		reg_103f4835_u0=1'h0;
reg		reg_6d11391e_u0=1'h0;
reg		reg_7a591648_u0=1'h0;
reg		reg_774d2b58_u0=1'h0;
reg		reg_32301a2a_u0=1'h0;
reg		reg_5cbbf0a1_u0=1'h0;
reg		reg_216d1570_u0=1'h0;
reg		reg_3e0fda11_u0=1'h0;
reg		reg_5e49be57_u0=1'h0;
reg		reg_09fdcdde_u0=1'h0;
reg		reg_62251200_u0=1'h0;
reg		reg_1e307217_u0=1'h0;
reg		reg_728582a2_u0=1'h0;
reg		reg_6bb9ab9e_u0=1'h0;
reg		reg_55d7a1ff_u0=1'h0;
reg		reg_2eee6ac6_u0=1'h0;
reg		reg_44cb88e0_u0=1'h0;
reg		reg_319759b9_u0=1'h0;
reg		reg_4bfc6bcc_u0=1'h0;
reg		reg_0dcebdfe_u0=1'h0;
reg		reg_08701441_u0=1'h0;
reg		reg_7a230a1a_u0=1'h0;
reg		reg_559271a8_u0=1'h0;
reg		reg_03167f2b_u0=1'h0;
reg		reg_0ffd27c0_u0=1'h0;
reg		reg_3711172f_u0=1'h0;
reg		reg_1340a77e_u0=1'h0;
reg		reg_7d9631d6_u0=1'h0;
reg		reg_69761137_u0=1'h0;
reg		reg_16db469f_u0=1'h0;
reg		reg_04257c62_u0=1'h0;
reg		reg_4cdea096_u0=1'h0;
reg		reg_6977313b_u0=1'h0;
reg		reg_297e0532_u0=1'h0;
reg		reg_54f5c8b9_u0=1'h0;
reg		reg_4db5d9f8_u0=1'h0;
reg		reg_188534c8_u0=1'h0;
reg		reg_32797234_u0=1'h0;
reg		reg_1fa5dbf4_u0=1'h0;
reg		reg_771e534d_u0=1'h0;
reg		reg_03167f2b_result_delayed_u0=1'h0;
reg		reg_1eb746e3_u0=1'h0;
reg		reg_2eee6ac6_result_delayed_u0=1'h0;
reg		reg_45429118_u0=1'h0;
reg		reg_1afd62a7_u0=1'h0;
reg		reg_0629ba72_u0=1'h0;
reg		reg_73b33bd3_u0=1'h0;
reg		reg_2159053d_u0=1'h0;
reg		reg_6da911c6_u0=1'h0;
reg		reg_1cdc40ac_u0=1'h0;
reg		reg_10ae20df_u0=1'h0;
reg		reg_41757d04_u0=1'h0;
reg		reg_306c2418_u0=1'h0;
reg		reg_5c0a547e_u0=1'h0;
reg		reg_20599c2d_u0=1'h0;
reg		reg_2586ddf0_u0=1'h0;
reg		reg_41757d04_result_delayed_u0=1'h0;
reg		reg_79dd91a5_u0=1'h0;
reg		reg_635d5720_u0=1'h0;
reg		reg_507b6cf9_u0=1'h0;
reg		reg_1340a77e_result_delayed_u0=1'h0;
reg		reg_04042082_u0=1'h0;
reg		reg_7080240a_u0=1'h0;
reg		reg_4cd5885f_u0=1'h0;
reg		reg_7080240a_result_delayed_u0=1'h0;
reg		reg_772bbfa5_u0=1'h0;
reg		reg_0dc8a158_u0=1'h0;
reg		reg_27cdb75f_u0=1'h0;
reg		reg_0e249eb7_u0=1'h0;
reg		reg_02d9964d_u0=1'h0;
reg		reg_50e04075_u0=1'h0;
reg		reg_33bcd31f_u0=1'h0;
reg		reg_19f2d151_u0=1'h0;
reg		reg_655155f8_u0=1'h0;
reg		reg_7432549f_u0=1'h0;
reg		reg_510951b8_u0=1'h0;
reg		reg_6ff27b40_u0=1'h0;
reg		reg_7bb0f302_u0=1'h0;
reg		reg_170037b2_u0=1'h0;
reg		reg_213ddd8e_u0=1'h0;
reg		reg_3d3f818b_u0=1'h0;
reg		reg_6f6443d2_u0=1'h0;
reg		reg_31278190_u0=1'h0;
reg		reg_4939b9f8_u0=1'h0;
reg		reg_73231fe1_u0=1'h0;
reg		reg_4cd5885f_result_delayed_u0=1'h0;
reg		reg_626c9aa9_u0=1'h0;
reg		reg_22e2922b_u0=1'h0;
reg		reg_5367bbad_u0=1'h0;
reg		reg_7368e3a4_u0=1'h0;
reg		reg_2e3a4ef5_u0=1'h0;
reg		reg_43dfbb10_u0=1'h0;
reg		reg_7d1e0dcf_u0=1'h0;
reg		reg_4ce52437_u0=1'h0;
reg		reg_745e0c57_result_delayed_u0=1'h0;
reg		reg_27394bed_u0=1'h0;
reg		reg_26de4e0b_u0=1'h0;
reg		reg_7b860f51_u0=1'h0;
reg		reg_1cdc40ac_result_delayed_u0=1'h0;
reg		reg_23b89b62_u0=1'h0;
reg		reg_3d75c9ae_u0=1'h0;
reg		reg_04042082_result_delayed_u0=1'h0;
reg		reg_49eb7136_u0=1'h0;
reg		reg_07979748_u0=1'h0;
reg		reg_561bf6ff_u0=1'h0;
reg		reg_32797234_result_delayed_u0=1'h0;
reg		reg_30e53c09_u0=1'h0;
reg		reg_01f9b917_u0=1'h0;
reg		reg_216d1570_result_delayed_u0=1'h0;
reg		reg_723816cc_u0=1'h0;
reg		reg_4bfc6bcc_result_delayed_u0=1'h0;
reg		reg_02179ae1_u0=1'h0;
reg		reg_608e408d_result_delayed_u0=1'h0;
reg		reg_2e3a4ef5_result_delayed_u0=1'h0;
reg		reg_5560159c_u0=1'h0;
reg		reg_776a1f94_u0=1'h0;
reg		reg_5c0a547e_result_delayed_u0=1'h0;
reg		reg_0da90157_u0=1'h0;
reg		reg_55d7a1ff_result_delayed_u0=1'h0;
reg		reg_2586ddf0_result_delayed_u0=1'h0;
reg		reg_619a949e_u0=1'h0;
reg		reg_414b944f_u0=1'h0;
reg		reg_00c68dc2_u0=1'h0;
reg		reg_13816284_u0=1'h0;
reg		reg_745e0c57_result_delayed_result_delayed_u0=1'h0;
reg		reg_10ae20df_result_delayed_u0=1'h0;
reg		reg_11b5ecb3_u0=1'h0;
reg		reg_662ef329_u0=1'h0;
reg		reg_56d52bdd_u0=1'h0;
reg		reg_11b5ecb3_result_delayed_u0=1'h0;
reg		reg_72f7e7fe_u0=1'h0;
reg		reg_7c98e992_u0=1'h0;
reg		reg_6f9f0292_u0=1'h0;
reg		reg_30251d3f_u0=1'h0;
reg		reg_4fd02acb_u0=1'h0;
reg		reg_1204a325_u0=1'h0;
reg		reg_6ccfd5e8_u0=1'h0;
reg		reg_0cc3a9eb_u0=1'h0;
reg		reg_63d04af9_u0=1'h0;
reg		reg_52cc27e6_u0=1'h0;
reg		reg_7107d82c_u0=1'h0;
reg		reg_32301a2a_result_delayed_u0=1'h0;
reg		reg_27e33acd_u0=1'h0;
reg		reg_56dbf3e8_u0=1'h0;
wire		or_u481_u0;
reg		reg_462c8f1b_u0=1'h0;
reg		reg_1340a77e_result_delayed_result_delayed_u0=1'h0;
reg		reg_7d792c42_u0=1'h0;
reg		reg_3711172f_result_delayed_u0=1'h0;
reg		reg_32797234_result_delayed_result_delayed_u0=1'h0;
reg		reg_10ff65be_u0=1'h0;
reg		reg_4d69442a_u0=1'h0;
reg		reg_6ca7ede4_u0=1'h0;
reg		reg_34313572_u0=1'h0;
reg		reg_328d47c8_u0=1'h0;
reg		reg_3bf5fabd_u0=1'h0;
reg		reg_27394bed_result_delayed_u0=1'h0;
reg		reg_107de137_u0=1'h0;
reg		reg_7a0a4746_u0=1'h0;
reg		reg_561bf6ff_result_delayed_u0=1'h0;
reg		reg_58245975_u0=1'h0;
reg		reg_2913cc47_u0=1'h0;
reg		reg_41757d04_result_delayed_result_delayed_u0=1'h0;
reg		reg_27cdb75f_result_delayed_u0=1'h0;
reg		reg_107de137_result_delayed_u0=1'h0;
reg		reg_0ffd27c0_result_delayed_u0=1'h0;
reg		reg_44a091fd_u0=1'h0;
reg		reg_30bea5e3_u0=1'h0;
reg		reg_2fe8a6b5_u0=1'h0;
reg		reg_55d7a1ff_result_delayed_result_delayed_u0=1'h0;
reg		reg_3ac9d797_u0=1'h0;
reg		reg_635d5720_result_delayed_u0=1'h0;
reg		reg_2913cc47_result_delayed_u0=1'h0;
reg		reg_306c2418_result_delayed_u0=1'h0;
reg		reg_4e506b37_u0=1'h0;
reg		reg_27faaa92_u0=1'h0;
reg		reg_107de137_result_delayed_result_delayed_u0=1'h0;
reg		reg_31f84093_u0=1'h0;
reg		reg_247a1111_u0=1'h0;
reg		reg_2fe8a6b5_result_delayed_u0=1'h0;
reg		reg_4a382354_u0=1'h0;
reg		reg_6b0d2e60_u0=1'h0;
reg		reg_5cbbf0a1_result_delayed_u0=1'h0;
reg		reg_7a0a4746_result_delayed_u0=1'h0;
reg		reg_619a949e_result_delayed_u0=1'h0;
reg		reg_5d3a8c49_u0=1'h0;
reg		reg_3d110516_result_delayed_u0=1'h0;
reg		reg_35c048b4_u0=1'h0;
reg		reg_49eb7136_result_delayed_u0=1'h0;
reg		reg_213ddd8e_result_delayed_u0=1'h0;
reg		reg_7c5e9123_u0=1'h0;
reg		reg_4692efed_u0=1'h0;
reg		reg_166d6bed_u0=1'h0;
reg		reg_47d1d653_u0=1'h0;
reg		reg_13e88a6a_u0=1'h0;
reg		reg_79dd91a5_result_delayed_u0=1'h0;
reg		reg_14ebcd6f_u0=1'h0;
reg		reg_157eb4fb_u0=1'h0;
reg		reg_32992b13_u0=1'h0;
reg		reg_1e3be3b6_u0=1'h0;
reg		reg_7ec5534b_u0=1'h0;
reg		reg_0d8e6001_u0=1'h0;
reg		reg_4cd5885f_result_delayed_result_delayed_u0=1'h0;
reg		reg_03bb9a29_u0=1'h0;
reg		reg_50412dd3_u0=1'h0;
reg		reg_322587b0_u0=1'h0;
reg		reg_3a122388_u0=1'h0;
reg		reg_1f4a72d1_u0=1'h0;
reg		reg_398e1010_u0=1'h0;
reg		reg_4bda7e7a_u0=1'h0;
reg		reg_6b0d2e60_result_delayed_u0=1'h0;
reg		reg_4b2b9289_u0=1'h0;
reg		reg_40236581_u0=1'h0;
reg		reg_7203dba7_u0=1'h0;
reg		reg_507b6cf9_result_delayed_u0=1'h0;
reg		reg_6e4f17e9_u0=1'h0;
reg		reg_12e5bf43_u0=1'h0;
reg		reg_4f83ce24_u0=1'h0;
reg		reg_774d2b58_result_delayed_u0=1'h0;
reg		reg_01f9b917_result_delayed_u0=1'h0;
reg		reg_776a1f94_result_delayed_u0=1'h0;
reg		reg_490168aa_u0=1'h0;
reg		reg_4bda7e7a_result_delayed_u0=1'h0;
reg		reg_5c0a547e_result_delayed_result_delayed_u0=1'h0;
reg		reg_6cdc1173_u0=1'h0;
reg		reg_5367bbad_result_delayed_u0=1'h0;
reg		reg_3365b2d6_u0=1'h0;
reg		reg_78922926_u0=1'h0;
reg		reg_4a747bcd_u0=1'h0;
reg		reg_37c4aa7f_u0=1'h0;
reg		reg_73231fe1_result_delayed_u0=1'h0;
reg		reg_33bcd31f_result_delayed_u0=1'h0;
reg		reg_1ba8b669_u0=1'h0;
reg		reg_4fd02acb_result_delayed_u0=1'h0;
reg		reg_35bbb476_u0=1'h0;
reg		reg_720d5fdc_u0=1'h0;
reg		reg_0f95e647_u0=1'h0;
reg		reg_5d1c80c9_u0=1'h0;
reg		reg_63d04af9_result_delayed_u0=1'h0;
reg		reg_2b4cee92_u0=1'h0;
reg		reg_20599c2d_result_delayed_u0=1'h0;
reg		reg_5c6cbd8d_u0=1'h0;
reg		reg_07979748_result_delayed_u0=1'h0;
reg		reg_7368e3a4_result_delayed_u0=1'h0;
reg		reg_1fa5dbf4_result_delayed_u0=1'h0;
reg		reg_1bd6ae3f_u0=1'h0;
reg		reg_4bf77a1c_u0=1'h0;
reg		reg_771e534d_result_delayed_u0=1'h0;
reg		reg_25c1902c_u0=1'h0;
reg		reg_68fe950f_u0=1'h0;
reg		reg_7984ac77_u0=1'h0;
reg		reg_32797234_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_7b860f51_result_delayed_u0=1'h0;
reg		reg_58245975_result_delayed_u0=1'h0;
reg		reg_626c9aa9_result_delayed_u0=1'h0;
reg		reg_728582a2_result_delayed_u0=1'h0;
reg		reg_04257c62_result_delayed_u0=1'h0;
reg		reg_4262839e_u0=1'h0;
reg		reg_74845d78_u0=1'h0;
reg		reg_248ca170_u0=1'h0;
reg		reg_0dcebdfe_result_delayed_u0=1'h0;
reg		reg_41757d04_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_2e9b949b_u0=1'h0;
reg		reg_739d919c_u0=1'h0;
reg		reg_12e5bf43_result_delayed_u0=1'h0;
reg		reg_0629ba72_result_delayed_u0=1'h0;
reg		reg_6da911c6_result_delayed_u0=1'h0;
reg		reg_43dfbb10_result_delayed_u0=1'h0;
reg		reg_776a1f94_result_delayed_result_delayed_u0=1'h0;
reg		reg_7a0a4746_result_delayed_result_delayed_u0=1'h0;
reg		reg_3771f97a_u0=1'h0;
reg		reg_248ca170_result_delayed_u0=1'h0;
reg		reg_5df5aff9_u0=1'h0;
reg		reg_5eb4b0ba_u0=1'h0;
reg		reg_2b82898d_u0=1'h0;
reg		reg_4692efed_result_delayed_u0=1'h0;
reg		reg_559271a8_result_delayed_u0=1'h0;
reg		reg_723816cc_result_delayed_u0=1'h0;
reg		reg_05d67bc0_u0=1'h0;
reg		reg_6ee280fb_u0=1'h0;
reg		reg_7a591648_result_delayed_u0=1'h0;
reg		reg_796d6b70_u0=1'h0;
reg		reg_6da911c6_result_delayed_result_delayed_u0=1'h0;
reg		reg_3562c342_u0=1'h0;
reg		reg_5cbbf0a1_result_delayed_result_delayed_u0=1'h0;
reg		reg_35875fa3_u0=1'h0;
reg		reg_328d47c8_result_delayed_u0=1'h0;
reg		reg_4cdea096_result_delayed_u0=1'h0;
reg		reg_103f4835_result_delayed_u0=1'h0;
reg		reg_1204a325_result_delayed_u0=1'h0;
reg		reg_64544e65_u0=1'h0;
reg		reg_655155f8_result_delayed_u0=1'h0;
reg		reg_31278190_result_delayed_u0=1'h0;
reg		reg_27410d75_u0=1'h0;
reg		reg_579fa5aa_u0=1'h0;
reg		reg_1e3be3b6_result_delayed_u0=1'h0;
reg		reg_02d9964d_result_delayed_u0=1'h0;
reg		reg_4db5d9f8_result_delayed_u0=1'h0;
reg		reg_3601783e_u0=1'h0;
reg		reg_08701441_result_delayed_u0=1'h0;
reg		reg_066f602e_u0=1'h0;
reg		reg_19f2d151_result_delayed_u0=1'h0;
reg		reg_7c98e992_result_delayed_u0=1'h0;
reg		reg_7c9a16d9_u0=1'h0;
reg		reg_343bd27c_u0=1'h0;
reg		reg_2b1f6158_u0=1'h0;
reg		reg_3c50f618_u0=1'h0;
reg		reg_3bf5fabd_result_delayed_u0=1'h0;
reg		reg_7c5e9123_result_delayed_u0=1'h0;
reg		reg_156fe33d_u0=1'h0;
reg		reg_4cdea096_result_delayed_result_delayed_u0=1'h0;
reg		reg_14ebcd6f_result_delayed_u0=1'h0;
reg		reg_170037b2_result_delayed_u0=1'h0;
reg		reg_30e53c09_result_delayed_u0=1'h0;
reg		reg_6fa9d1fe_u0=1'h0;
reg		reg_36d51882_u0=1'h0;
reg		reg_4262839e_result_delayed_u0=1'h0;
reg		reg_65390362_u0=1'h0;
reg		reg_00c68dc2_result_delayed_u0=1'h0;
reg		reg_6f9f0292_result_delayed_u0=1'h0;
reg		reg_2711b972_u0=1'h0;
reg		reg_33bcd31f_result_delayed_result_delayed_u0=1'h0;
reg		reg_2eee6ac6_result_delayed_result_delayed_u0=1'h0;
reg		reg_357d771a_u0=1'h0;
reg		reg_5bf74d9f_u0=1'h0;
reg		reg_0ba46dcc_u0=1'h0;
reg		reg_7d792c42_result_delayed_u0=1'h0;
reg		reg_772bbfa5_result_delayed_u0=1'h0;
reg		reg_1d5ae331_u0=1'h0;
reg		reg_0da887c4_u0=1'h0;
reg		reg_32301a2a_result_delayed_result_delayed_u0=1'h0;
reg		reg_41a8efc6_u0=1'h0;
reg		reg_7bb0f302_result_delayed_u0=1'h0;
reg		reg_6bb9ab9e_result_delayed_u0=1'h0;
reg		reg_71343346_u0=1'h0;
reg		reg_2f9c95e8_u0=1'h0;
reg		reg_0178db0e_u0=1'h0;
reg		reg_5eb4b0ba_result_delayed_u0=1'h0;
reg		reg_02d9964d_result_delayed_result_delayed_u0=1'h0;
reg		reg_27394bed_result_delayed_result_delayed_u0=1'h0;
reg		reg_68fe950f_result_delayed_u0=1'h0;
reg		reg_7bb0f302_result_delayed_result_delayed_u0=1'h0;
reg		reg_45429118_result_delayed_u0=1'h0;
reg		reg_19f2d151_result_delayed_result_delayed_u0=1'h0;
reg		reg_32992b13_result_delayed_u0=1'h0;
reg		reg_10ae20df_result_delayed_result_delayed_u0=1'h0;
reg		reg_1e3be3b6_result_delayed_result_delayed_u0=1'h0;
reg		reg_56d52bdd_result_delayed_u0=1'h0;
reg		reg_6b0d2e60_result_delayed_result_delayed_u0=1'h0;
reg		reg_7a230a1a_result_delayed_u0=1'h0;
reg		reg_0ba46dcc_result_delayed_u0=1'h0;
reg		reg_247e36e9_u0=1'h0;
reg		reg_248ca170_result_delayed_result_delayed_u0=1'h0;
reg		reg_43dfbb10_result_delayed_result_delayed_u0=1'h0;
reg		reg_490168aa_result_delayed_u0=1'h0;
reg		reg_4cd5885f_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_4262839e_result_delayed_result_delayed_u0=1'h0;
reg		reg_31f84093_result_delayed_u0=1'h0;
reg		reg_3d3b97a5_u0=1'h0;
reg		reg_02179ae1_result_delayed_u0=1'h0;
reg		reg_561bf6ff_result_delayed_result_delayed_u0=1'h0;
reg		reg_03167f2b_result_delayed_result_delayed_u0=1'h0;
reg		reg_4ce52437_result_delayed_u0=1'h0;
reg		reg_19f2d151_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_6ca7ede4_result_delayed_u0=1'h0;
reg		reg_0ef60446_u0=1'h0;
reg		reg_2fe8a6b5_result_delayed_result_delayed_u0=1'h0;
reg		reg_6ff27b40_result_delayed_u0=1'h0;
reg		reg_4cdea096_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_5cbbf0a1_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_7432549f_result_delayed_u0=1'h0;
reg		reg_6ee42c26_u0=1'h0;
reg		reg_4692efed_result_delayed_result_delayed_u0=1'h0;
reg		reg_0c928251_u0=1'h0;
reg		reg_20599c2d_result_delayed_result_delayed_u0=1'h0;
reg		reg_319759b9_result_delayed_u0=1'h0;
reg		reg_62251200_result_delayed_u0=1'h0;
reg		reg_7d792c42_result_delayed_result_delayed_u0=1'h0;
reg		reg_1fa5dbf4_result_delayed_result_delayed_u0=1'h0;
reg		reg_5eb4b0ba_result_delayed_result_delayed_u0=1'h0;
reg		reg_3dfa0f2c_u0=1'h0;
reg		reg_55d7a1ff_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_6ee42c26_result_delayed_u0=1'h0;
reg		reg_26bc9067_u0=1'h0;
reg		reg_1ba8b669_result_delayed_u0=1'h0;
reg		reg_3d75c9ae_result_delayed_u0=1'h0;
reg		reg_31f84093_result_delayed_result_delayed_u0=1'h0;
reg		reg_42f3b02c_u0=1'h0;
reg		reg_2afa8c1b_u0=1'h0;
reg		reg_7c5e9123_result_delayed_result_delayed_u0=1'h0;
reg		reg_2ab2a055_u0=1'h0;
reg		reg_69761137_result_delayed_u0=1'h0;
reg		reg_561ae0f2_u0=1'h0;
reg		reg_1eb746e3_result_delayed_u0=1'h0;
reg		reg_10ff65be_result_delayed_u0=1'h0;
reg		reg_4e506b37_result_delayed_u0=1'h0;
reg		reg_3a122388_result_delayed_u0=1'h0;
reg		reg_31f84093_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_0ae85810_u0=1'h0;
reg		reg_3c50f618_result_delayed_u0=1'h0;
reg		reg_4692efed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_6f6443d2_result_delayed_u0=1'h0;
reg		reg_4d69442a_result_delayed_u0=1'h0;
reg		reg_3cd29fd9_u0=1'h0;
reg		reg_73b33bd3_result_delayed_u0=1'h0;
reg		reg_25c1902c_result_delayed_u0=1'h0;
reg		reg_729e0d87_u0=1'h0;
reg		reg_30bea5e3_result_delayed_u0=1'h0;
reg		reg_44cb88e0_result_delayed_u0=1'h0;
reg		reg_606de772_u0=1'h0;
wire		and_u1764_u0;
reg		reg_71343346_result_delayed_u0=1'h0;
reg		reg_49eb7136_result_delayed_result_delayed_u0=1'h0;
reg		reg_2586ddf0_result_delayed_result_delayed_u0=1'h0;
reg		reg_7352b877_u0=1'h0;
reg		reg_40236581_result_delayed_u0=1'h0;
reg		reg_414b944f_result_delayed_u0=1'h0;
reg		reg_739d919c_result_delayed_u0=1'h0;
reg		reg_3cd29fd9_result_delayed_u0=1'h0;
reg		reg_188534c8_result_delayed_u0=1'h0;
reg		reg_09fdcdde_result_delayed_u0=1'h0;
reg		reg_43d7d4e5_u0=1'h0;
reg		reg_02179ae1_result_delayed_result_delayed_u0=1'h0;
wire		mux_u180;
wire		or_u482_u0;
reg		reg_22387d0e_u0=1'h0;
reg		reg_32301a2a_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_357d771a_result_delayed_u0=1'h0;
reg		reg_5e49be57_result_delayed_u0=1'h0;
reg		reg_776a1f94_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_552e2e6e_u0=1'h0;
reg		reg_2711b972_result_delayed_u0=1'h0;
reg		reg_398e1010_result_delayed_u0=1'h0;
reg		reg_78922926_result_delayed_u0=1'h0;
reg		reg_630a4c43_u0=1'h0;
reg		reg_4939b9f8_result_delayed_u0=1'h0;
reg		reg_0da90157_result_delayed_u0=1'h0;
reg		reg_635d5720_result_delayed_result_delayed_u0=1'h0;
reg		reg_343bd27c_result_delayed_u0=1'h0;
reg		reg_3e0fda11_result_delayed_u0=1'h0;
reg		reg_3ac9d797_result_delayed_u0=1'h0;
reg		reg_3d3b97a5_result_delayed_u0=1'h0;
reg		reg_3562c342_result_delayed_u0=1'h0;
reg		reg_157eb4fb_result_delayed_u0=1'h0;
reg		reg_6ccfd5e8_result_delayed_u0=1'h0;
reg		reg_2b2ea879_u0=1'h0;
reg		reg_02179ae1_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_626c9aa9_result_delayed_result_delayed_u0=1'h0;
reg		reg_4e506b37_result_delayed_result_delayed_u0=1'h0;
reg		reg_2159053d_result_delayed_u0=1'h0;
reg		reg_7ec5534b_result_delayed_u0=1'h0;
reg		reg_0ffd27c0_result_delayed_result_delayed_u0=1'h0;
reg		reg_32797234_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_3d110516_result_delayed_result_delayed_u0=1'h0;
reg		reg_7080240a_result_delayed_result_delayed_u0=1'h0;
reg		reg_55d7a1ff_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_6ca7ede4_result_delayed_result_delayed_u0=1'h0;
reg		reg_23b89b62_result_delayed_u0=1'h0;
reg		reg_1afd62a7_result_delayed_u0=1'h0;
reg		reg_35875fa3_result_delayed_u0=1'h0;
reg		reg_579fa5aa_result_delayed_u0=1'h0;
reg		reg_2e3a4ef5_result_delayed_result_delayed_u0=1'h0;
reg		reg_772bbfa5_result_delayed_result_delayed_u0=1'h0;
reg		reg_50e04075_result_delayed_u0=1'h0;
reg		reg_1bd6ae3f_result_delayed_u0=1'h0;
reg		reg_326d6def_u0=1'h0;
reg		reg_6e4f17e9_result_delayed_u0=1'h0;
reg		reg_608e408d_result_delayed_result_delayed_u0=1'h0;
reg		reg_7d792c42_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_066f602e_result_delayed_u0=1'h0;
reg		reg_2a9c2111_u0=1'h0;
reg		reg_248ca170_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_6da911c6_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_4bc0004f_u0=1'h0;
reg		reg_04257c62_result_delayed_result_delayed_u0=1'h0;
reg		reg_3a122388_result_delayed_result_delayed_u0=1'h0;
reg		reg_056e42f2_u0=1'h0;
reg		reg_319759b9_result_delayed_result_delayed_u0=1'h0;
reg		reg_4db5d9f8_result_delayed_result_delayed_u0=1'h0;
reg		reg_510951b8_result_delayed_u0=1'h0;
reg		reg_22e2922b_result_delayed_u0=1'h0;
reg		reg_6d11391e_result_delayed_u0=1'h0;
reg		reg_1e307217_result_delayed_u0=1'h0;
reg		reg_2b82898d_result_delayed_u0=1'h0;
reg		reg_1d5ae331_result_delayed_u0=1'h0;
reg		reg_41757d04_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_157eb4fb_result_delayed_result_delayed_u0=1'h0;
reg		reg_4a382354_result_delayed_u0=1'h0;
wire		and_u1765_u0;
reg		reg_0e249eb7_result_delayed_u0=1'h0;
reg		reg_1bd6ae3f_result_delayed_result_delayed_u0=1'h0;
reg		reg_2c6d2fd0_u0=1'h0;
reg		reg_0dc8a158_result_delayed_u0=1'h0;
reg		reg_216d1570_result_delayed_result_delayed_u0=1'h0;
reg		reg_72f7e7fe_result_delayed_u0=1'h0;
reg		reg_2ab2a055_result_delayed_u0=1'h0;
reg		reg_2b4cee92_result_delayed_u0=1'h0;
reg		reg_16db469f_result_delayed_u0=1'h0;
reg		reg_4bc0004f_result_delayed_u0=1'h0;
reg		reg_2e9b949b_result_delayed_u0=1'h0;
reg		reg_07979748_result_delayed_result_delayed_u0=1'h0;
reg		reg_4bfc6bcc_result_delayed_result_delayed_u0=1'h0;
reg		reg_297e0532_result_delayed_u0=1'h0;
reg		reg_1bd6ae3f_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_776a1f94_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_74845d78_result_delayed_u0=1'h0;
reg		reg_247a1111_result_delayed_u0=1'h0;
reg		reg_30bea5e3_result_delayed_result_delayed_u0=1'h0;
reg		reg_170037b2_result_delayed_result_delayed_u0=1'h0;
reg		reg_319759b9_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_63d04af9_result_delayed_result_delayed_u0=1'h0;
reg		reg_6ee280fb_result_delayed_u0=1'h0;
reg		reg_3771f97a_result_delayed_u0=1'h0;
reg		reg_44a091fd_result_delayed_u0=1'h0;
reg		reg_5c0a547e_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_7a591648_result_delayed_result_delayed_u0=1'h0;
wire		or_u483_u0;
wire		or_u484_u0;
wire		mux_u181_u0;
wire		or_u485_u0;
wire		and_u1766_u0;
reg		and_delayed_u118=1'h0;
reg		and_delayed_result_delayed_u9=1'h0;
wire		and_u1767_u0;
wire		or_u486_u0;
wire	[31:0]	mux_u182_u0;
wire		or_u487_u0;
reg		and_delayed_result_delayed_result_delayed_u2=1'h0;
wire		or_u488_u0;
wire		and_u1768_u0;
wire		or_u489_u0;
reg		and_delayed_u119_u0=1'h0;
wire		and_u1769_u0;
wire signed	[31:0]	equals_u94_a_signed;
wire signed	[31:0]	equals_u94_b_signed;
wire		equals_u94;
wire		and_u1770_u0;
wire		and_u1771_u0;
wire		not_u350_u0;
wire		and_u1772_u0;
wire		and_u1773_u0;
wire		not_u351_u0;
wire		lessThan_u39;
wire signed	[31:0]	lessThan_u39_a_signed;
wire signed	[31:0]	lessThan_u39_b_signed;
wire		not_u352_u0;
wire		and_u1774_u0;
wire		and_u1775_u0;
wire		not_u353_u0;
wire		and_u1776_u0;
wire		and_u1777_u0;
wire	[31:0]	add;
wire		and_u1778_u0;
wire	[15:0]	simplePinWrite_u318;
wire	[15:0]	simplePinWrite_u319;
wire		simplePinWrite_u320;
wire	[31:0]	add_u68;
reg	[15:0]	syncEnable_u180=16'h0;
wire	[15:0]	mux_u183_u0;
wire		and_u1779_u0;
wire		and_u1780_u0;
reg	[15:0]	syncEnable_u181_u0=16'h0;
reg		and_delayed_u120_u0=1'h0;
reg		and_delayed_u121_u0=1'h0;
reg	[31:0]	syncEnable_u182_u0=32'h0;
wire	[15:0]	mux_u184_u0;
reg		reg_4dcef723_u0=1'h0;
reg		reg_645b9fd5_u0=1'h0;
wire		and_u1781_u0;
reg	[15:0]	syncEnable_u183_u0=16'h0;
wire		and_u1782_u0;
wire	[31:0]	mux_u185_u0;
reg		reg_1a01de45_u0=1'h0;
reg		reg_535070be_u0=1'h0;
reg	[31:0]	syncEnable_u184_u0=32'h0;
wire		and_u1783_u0;
wire		and_u1784_u0;
wire	[31:0]	mux_u186_u0;
wire	[15:0]	mux_u187_u0;
reg	[15:0]	syncEnable_u185_u0=16'h0;
wire	[15:0]	mux_u188_u0;
reg		reg_5039c73f_u0=1'h0;
wire		and_u1785_u0;
reg	[31:0]	syncEnable_u186_u0=32'h0;
wire		and_u1786_u0;
wire	[31:0]	mux_u189_u0;
reg		and_delayed_u122_u0=1'h0;
reg	[15:0]	syncEnable_u187_u0=16'h0;
wire		mux_u190_u0;
wire		or_u490_u0;
wire	[15:0]	latch_4d9bcb18_out;
reg	[15:0]	latch_4d9bcb18_reg=16'h0;
wire		or_u491_u0;
wire	[31:0]	mux_u191_u0;
wire	[31:0]	latch_1e7607d8_out;
reg	[31:0]	latch_1e7607d8_reg=32'h0;
wire		or_u492_u0;
wire		mux_u192_u0;
reg		block_GO_delayed_u6=1'h0;
wire		or_u493_u0;
wire	[31:0]	mux_u193_u0;
wire	[31:0]	mux_u194_u0;
wire		or_u494_u0;
reg	[31:0]	fbReg_temp_fsmOldState_resized_HH1_xy_3_u0=32'h0;
reg		loopControl_u3=1'h0;
wire	[15:0]	mux_u195_u0;
reg		syncEnable_u188_u0=1'h0;
reg	[15:0]	fbReg_Out1Portvalue_u0=16'h0;
reg		reg_36b6d836_u0=1'h0;
wire		or_u495_u0;
wire	[31:0]	mux_u196_u0;
wire		or_u496_u0;
reg		reg_36b6d836_result_delayed_u0=1'h0;
wire		or_u497_u0;
wire	[31:0]	mux_u197_u0;
wire		or_u498_u0;
wire		mux_u198_u0;
wire		or_u499_u0;
wire		mux_u199_u0;
assign and_u1754_u0=or_u494_u0&or_u494_u0;
assign lessThan_a_unsigned=port_0fbd4927_;
assign lessThan_b_unsigned=16'h100;
assign lessThan=lessThan_a_unsigned<lessThan_b_unsigned;
assign equals_a_unsigned=port_0fbd4927_;
assign equals_b_unsigned=16'h100;
assign equals=equals_a_unsigned==equals_b_unsigned;
assign lessThan_u38_a_unsigned=port_0d76a61b_;
assign lessThan_u38_b_unsigned=16'h2;
assign lessThan_u38=lessThan_u38_a_unsigned<lessThan_u38_b_unsigned;
assign andOp=equals&lessThan_u38;
assign equals_u92_a_unsigned=port_0d76a61b_;
assign equals_u92_b_unsigned=16'h2;
assign equals_u92=equals_u92_a_unsigned==equals_u92_b_unsigned;
assign equals_u93_a_signed={31'b0, port_0712fa18_};
assign equals_u93_b_signed=32'h0;
assign equals_u93=equals_u93_a_signed==equals_u93_b_signed;
assign not_u346_u0=~equals_u93;
assign and_u1755_u0=and_u1754_u0&equals_u93;
assign and_u1756_u0=and_u1754_u0&not_u346_u0;
assign andOp_u113=lessThan&port_316bbc7c_;
assign not_u347_u0=~andOp_u113;
assign and_u1757_u0=and_u1769_u0&not_u347_u0;
assign and_u1758_u0=and_u1769_u0&andOp_u113;
assign simplePinWrite=and_u1766_u0&{1{and_u1766_u0}};
assign and_u1759_u0=and_u1767_u0&andOp;
assign and_u1760_u0=and_u1767_u0&not_u348_u0;
assign not_u348_u0=~andOp;
assign simplePinWrite_u316=and_u1765_u0&{1{and_u1765_u0}};
assign and_u1761_u0=and_u1764_u0&equals_u92;
assign not_u349_u0=~equals_u92;
assign and_u1762_u0=and_u1764_u0&not_u349_u0;
assign simplePinWrite_u317=and_u1763_u0&{1{and_u1763_u0}};
assign and_u1763_u0=and_u1761_u0&and_u1764_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_608e408d_u0<=1'h0;
else reg_608e408d_u0<=reg_6f6443d2_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3d110516_u0<=1'h0;
else reg_3d110516_u0<=reg_54f5c8b9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_745e0c57_u0<=1'h0;
else reg_745e0c57_u0<=reg_32301a2a_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_103f4835_u0<=1'h0;
else reg_103f4835_u0<=reg_4f83ce24_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6d11391e_u0<=1'h0;
else reg_6d11391e_u0<=reg_26de4e0b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a591648_u0<=1'h0;
else reg_7a591648_u0<=reg_12e5bf43_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_774d2b58_u0<=1'h0;
else reg_774d2b58_u0<=reg_107de137_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_32301a2a_u0<=1'h0;
else reg_32301a2a_u0<=reg_1cdc40ac_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5cbbf0a1_u0<=1'h0;
else reg_5cbbf0a1_u0<=reg_11b5ecb3_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_216d1570_u0<=1'h0;
else reg_216d1570_u0<=reg_13816284_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3e0fda11_u0<=1'h0;
else reg_3e0fda11_u0<=reg_47d1d653_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5e49be57_u0<=1'h0;
else reg_5e49be57_u0<=reg_745e0c57_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_09fdcdde_u0<=1'h0;
else reg_09fdcdde_u0<=reg_7d9631d6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_62251200_u0<=1'h0;
else reg_62251200_u0<=reg_606de772_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1e307217_u0<=1'h0;
else reg_1e307217_u0<=reg_626c9aa9_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_728582a2_u0<=1'h0;
else reg_728582a2_u0<=reg_2913cc47_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6bb9ab9e_u0<=1'h0;
else reg_6bb9ab9e_u0<=reg_27cdb75f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_55d7a1ff_u0<=1'h0;
else reg_55d7a1ff_u0<=reg_729e0d87_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2eee6ac6_u0<=1'h0;
else reg_2eee6ac6_u0<=reg_2b2ea879_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_44cb88e0_u0<=1'h0;
else reg_44cb88e0_u0<=reg_2ab2a055_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_319759b9_u0<=1'h0;
else reg_319759b9_u0<=reg_30e53c09_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4bfc6bcc_u0<=1'h0;
else reg_4bfc6bcc_u0<=reg_50412dd3_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0dcebdfe_u0<=1'h0;
else reg_0dcebdfe_u0<=reg_739d919c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_08701441_u0<=1'h0;
else reg_08701441_u0<=reg_62251200_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a230a1a_u0<=1'h0;
else reg_7a230a1a_u0<=reg_14ebcd6f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_559271a8_u0<=1'h0;
else reg_559271a8_u0<=reg_247e36e9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_03167f2b_u0<=1'h0;
else reg_03167f2b_u0<=reg_5bf74d9f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0ffd27c0_u0<=1'h0;
else reg_0ffd27c0_u0<=reg_3562c342_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3711172f_u0<=1'h0;
else reg_3711172f_u0<=reg_04042082_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1340a77e_u0<=1'h0;
else reg_1340a77e_u0<=reg_328d47c8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7d9631d6_u0<=1'h0;
else reg_7d9631d6_u0<=reg_79dd91a5_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_69761137_u0<=1'h0;
else reg_69761137_u0<=reg_4d69442a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_16db469f_u0<=1'h0;
else reg_16db469f_u0<=reg_3e0fda11_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_04257c62_u0<=1'h0;
else reg_04257c62_u0<=reg_0d8e6001_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4cdea096_u0<=1'h0;
else reg_4cdea096_u0<=reg_6977313b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6977313b_u0<=1'h0;
else reg_6977313b_u0<=reg_2e9b949b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_297e0532_u0<=1'h0;
else reg_297e0532_u0<=reg_056e42f2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_54f5c8b9_u0<=1'h0;
else reg_54f5c8b9_u0<=reg_0dc8a158_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4db5d9f8_u0<=1'h0;
else reg_4db5d9f8_u0<=reg_35875fa3_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_188534c8_u0<=1'h0;
else reg_188534c8_u0<=reg_19f2d151_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_32797234_u0<=1'h0;
else reg_32797234_u0<=reg_490168aa_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1fa5dbf4_u0<=1'h0;
else reg_1fa5dbf4_u0<=reg_772bbfa5_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_771e534d_u0<=1'h0;
else reg_771e534d_u0<=reg_3711172f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_03167f2b_result_delayed_u0<=1'h0;
else reg_03167f2b_result_delayed_u0<=reg_03167f2b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1eb746e3_u0<=1'h0;
else reg_1eb746e3_u0<=reg_4db5d9f8_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2eee6ac6_result_delayed_u0<=1'h0;
else reg_2eee6ac6_result_delayed_u0<=reg_2eee6ac6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_45429118_u0<=1'h0;
else reg_45429118_u0<=reg_2afa8c1b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1afd62a7_u0<=1'h0;
else reg_1afd62a7_u0<=reg_10ff65be_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0629ba72_u0<=1'h0;
else reg_0629ba72_u0<=reg_5560159c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_73b33bd3_u0<=1'h0;
else reg_73b33bd3_u0<=reg_03bb9a29_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2159053d_u0<=1'h0;
else reg_2159053d_u0<=reg_27faaa92_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6da911c6_u0<=1'h0;
else reg_6da911c6_u0<=reg_188534c8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1cdc40ac_u0<=1'h0;
else reg_1cdc40ac_u0<=reg_41a8efc6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_10ae20df_u0<=1'h0;
else reg_10ae20df_u0<=reg_357d771a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_41757d04_u0<=1'h0;
else reg_41757d04_u0<=reg_20599c2d_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_306c2418_u0<=1'h0;
else reg_306c2418_u0<=reg_771e534d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5c0a547e_u0<=1'h0;
else reg_5c0a547e_u0<=reg_3d3f818b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_20599c2d_u0<=1'h0;
else reg_20599c2d_u0<=reg_1f4a72d1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2586ddf0_u0<=1'h0;
else reg_2586ddf0_u0<=reg_26bc9067_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_41757d04_result_delayed_u0<=1'h0;
else reg_41757d04_result_delayed_u0<=reg_41757d04_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_79dd91a5_u0<=1'h0;
else reg_79dd91a5_u0<=reg_0cc3a9eb_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_635d5720_u0<=1'h0;
else reg_635d5720_u0<=reg_34313572_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_507b6cf9_u0<=1'h0;
else reg_507b6cf9_u0<=reg_4939b9f8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1340a77e_result_delayed_u0<=1'h0;
else reg_1340a77e_result_delayed_u0<=reg_1340a77e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_04042082_u0<=1'h0;
else reg_04042082_u0<=reg_52cc27e6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7080240a_u0<=1'h0;
else reg_7080240a_u0<=reg_213ddd8e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4cd5885f_u0<=1'h0;
else reg_4cd5885f_u0<=reg_5c6cbd8d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7080240a_result_delayed_u0<=1'h0;
else reg_7080240a_result_delayed_u0<=reg_7080240a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_772bbfa5_u0<=1'h0;
else reg_772bbfa5_u0<=reg_7ec5534b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0dc8a158_u0<=1'h0;
else reg_0dc8a158_u0<=reg_662ef329_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_27cdb75f_u0<=1'h0;
else reg_27cdb75f_u0<=reg_0ffd27c0_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0e249eb7_u0<=1'h0;
else reg_0e249eb7_u0<=reg_13e88a6a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_02d9964d_u0<=1'h0;
else reg_02d9964d_u0<=reg_3d75c9ae_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_50e04075_u0<=1'h0;
else reg_50e04075_u0<=reg_30251d3f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_33bcd31f_u0<=1'h0;
else reg_33bcd31f_u0<=reg_1340a77e_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_19f2d151_u0<=1'h0;
else reg_19f2d151_u0<=reg_507b6cf9_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_655155f8_u0<=1'h0;
else reg_655155f8_u0<=reg_2e3a4ef5_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7432549f_u0<=1'h0;
else reg_7432549f_u0<=reg_7a230a1a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_510951b8_u0<=1'h0;
else reg_510951b8_u0<=reg_1ba8b669_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6ff27b40_u0<=1'h0;
else reg_6ff27b40_u0<=reg_68fe950f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7bb0f302_u0<=1'h0;
else reg_7bb0f302_u0<=reg_33bcd31f_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_170037b2_u0<=1'h0;
else reg_170037b2_u0<=reg_774d2b58_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_213ddd8e_u0<=1'h0;
else reg_213ddd8e_u0<=reg_462c8f1b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3d3f818b_u0<=1'h0;
else reg_3d3f818b_u0<=reg_322587b0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6f6443d2_u0<=1'h0;
else reg_6f6443d2_u0<=reg_58245975_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_31278190_u0<=1'h0;
else reg_31278190_u0<=reg_166d6bed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4939b9f8_u0<=1'h0;
else reg_4939b9f8_u0<=reg_1204a325_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_73231fe1_u0<=1'h0;
else reg_73231fe1_u0<=reg_7c9a16d9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4cd5885f_result_delayed_u0<=1'h0;
else reg_4cd5885f_result_delayed_u0<=reg_4cd5885f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_626c9aa9_u0<=1'h0;
else reg_626c9aa9_u0<=reg_44a091fd_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_22e2922b_u0<=1'h0;
else reg_22e2922b_u0<=reg_35c048b4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5367bbad_u0<=1'h0;
else reg_5367bbad_u0<=reg_32992b13_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7368e3a4_u0<=1'h0;
else reg_7368e3a4_u0<=reg_7d1e0dcf_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2e3a4ef5_u0<=1'h0;
else reg_2e3a4ef5_u0<=reg_45429118_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_43dfbb10_u0<=1'h0;
else reg_43dfbb10_u0<=reg_6cdc1173_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7d1e0dcf_u0<=1'h0;
else reg_7d1e0dcf_u0<=reg_6ff27b40_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4ce52437_u0<=1'h0;
else reg_4ce52437_u0<=reg_510951b8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_745e0c57_result_delayed_u0<=1'h0;
else reg_745e0c57_result_delayed_u0<=reg_745e0c57_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_27394bed_u0<=1'h0;
else reg_27394bed_u0<=reg_41757d04_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_26de4e0b_u0<=1'h0;
else reg_26de4e0b_u0<=reg_4ce52437_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7b860f51_u0<=1'h0;
else reg_7b860f51_u0<=reg_720d5fdc_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1cdc40ac_result_delayed_u0<=1'h0;
else reg_1cdc40ac_result_delayed_u0<=reg_1cdc40ac_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_23b89b62_u0<=1'h0;
else reg_23b89b62_u0<=reg_27e33acd_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3d75c9ae_u0<=1'h0;
else reg_3d75c9ae_u0<=reg_6fa9d1fe_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_04042082_result_delayed_u0<=1'h0;
else reg_04042082_result_delayed_u0<=reg_04042082_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_49eb7136_u0<=1'h0;
else reg_49eb7136_u0<=reg_398e1010_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_07979748_u0<=1'h0;
else reg_07979748_u0<=reg_066f602e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_561bf6ff_u0<=1'h0;
else reg_561bf6ff_u0<=reg_306c2418_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_32797234_result_delayed_u0<=1'h0;
else reg_32797234_result_delayed_u0<=reg_32797234_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_30e53c09_u0<=1'h0;
else reg_30e53c09_u0<=reg_35bbb476_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01f9b917_u0<=1'h0;
else reg_01f9b917_u0<=reg_0f95e647_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_216d1570_result_delayed_u0<=1'h0;
else reg_216d1570_result_delayed_u0<=reg_216d1570_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_723816cc_u0<=1'h0;
else reg_723816cc_u0<=reg_7c98e992_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4bfc6bcc_result_delayed_u0<=1'h0;
else reg_4bfc6bcc_result_delayed_u0<=reg_4bfc6bcc_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_02179ae1_u0<=1'h0;
else reg_02179ae1_u0<=reg_05d67bc0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_608e408d_result_delayed_u0<=1'h0;
else reg_608e408d_result_delayed_u0<=reg_608e408d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2e3a4ef5_result_delayed_u0<=1'h0;
else reg_2e3a4ef5_result_delayed_u0<=reg_2e3a4ef5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5560159c_u0<=1'h0;
else reg_5560159c_u0<=reg_2a9c2111_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_776a1f94_u0<=1'h0;
else reg_776a1f94_u0<=reg_0ae85810_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5c0a547e_result_delayed_u0<=1'h0;
else reg_5c0a547e_result_delayed_u0<=reg_5c0a547e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0da90157_u0<=1'h0;
else reg_0da90157_u0<=reg_7352b877_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_55d7a1ff_result_delayed_u0<=1'h0;
else reg_55d7a1ff_result_delayed_u0<=reg_55d7a1ff_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2586ddf0_result_delayed_u0<=1'h0;
else reg_2586ddf0_result_delayed_u0<=reg_2586ddf0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_619a949e_u0<=1'h0;
else reg_619a949e_u0<=reg_6b0d2e60_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_414b944f_u0<=1'h0;
else reg_414b944f_u0<=reg_56dbf3e8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00c68dc2_u0<=1'h0;
else reg_00c68dc2_u0<=reg_1bd6ae3f_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_13816284_u0<=1'h0;
else reg_13816284_u0<=reg_7107d82c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_745e0c57_result_delayed_result_delayed_u0<=1'h0;
else reg_745e0c57_result_delayed_result_delayed_u0<=reg_745e0c57_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_10ae20df_result_delayed_u0<=1'h0;
else reg_10ae20df_result_delayed_u0<=reg_10ae20df_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_11b5ecb3_u0<=1'h0;
else reg_11b5ecb3_u0<=reg_2711b972_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_662ef329_u0<=1'h0;
else reg_662ef329_u0<=reg_2f9c95e8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_56d52bdd_u0<=1'h0;
else reg_56d52bdd_u0<=reg_7d792c42_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_11b5ecb3_result_delayed_u0<=1'h0;
else reg_11b5ecb3_result_delayed_u0<=reg_11b5ecb3_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_72f7e7fe_u0<=1'h0;
else reg_72f7e7fe_u0<=reg_552e2e6e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7c98e992_u0<=1'h0;
else reg_7c98e992_u0<=reg_4fd02acb_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6f9f0292_u0<=1'h0;
else reg_6f9f0292_u0<=reg_170037b2_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_30251d3f_u0<=1'h0;
else reg_30251d3f_u0<=reg_1fa5dbf4_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4fd02acb_u0<=1'h0;
else reg_4fd02acb_u0<=reg_0629ba72_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1204a325_u0<=1'h0;
else reg_1204a325_u0<=reg_2b1f6158_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6ccfd5e8_u0<=1'h0;
else reg_6ccfd5e8_u0<=reg_4a382354_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0cc3a9eb_u0<=1'h0;
else reg_0cc3a9eb_u0<=reg_2b82898d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_63d04af9_u0<=1'h0;
else reg_63d04af9_u0<=reg_4bfc6bcc_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_52cc27e6_u0<=1'h0;
else reg_52cc27e6_u0<=reg_7203dba7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7107d82c_u0<=1'h0;
else reg_7107d82c_u0<=reg_630a4c43_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_32301a2a_result_delayed_u0<=1'h0;
else reg_32301a2a_result_delayed_u0<=reg_32301a2a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_27e33acd_u0<=1'h0;
else reg_27e33acd_u0<=reg_6ccfd5e8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_56dbf3e8_u0<=1'h0;
else reg_56dbf3e8_u0<=reg_6ca7ede4_result_delayed_result_delayed_u0;
end
assign or_u481_u0=reg_3365b2d6_u0|reg_27410d75_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_462c8f1b_u0<=1'h0;
else reg_462c8f1b_u0<=reg_5d1c80c9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1340a77e_result_delayed_result_delayed_u0<=1'h0;
else reg_1340a77e_result_delayed_result_delayed_u0<=reg_1340a77e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7d792c42_u0<=1'h0;
else reg_7d792c42_u0<=reg_4a747bcd_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3711172f_result_delayed_u0<=1'h0;
else reg_3711172f_result_delayed_u0<=reg_3711172f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_32797234_result_delayed_result_delayed_u0<=1'h0;
else reg_32797234_result_delayed_result_delayed_u0<=reg_32797234_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_10ff65be_u0<=1'h0;
else reg_10ff65be_u0<=reg_32797234_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4d69442a_u0<=1'h0;
else reg_4d69442a_u0<=reg_728582a2_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6ca7ede4_u0<=1'h0;
else reg_6ca7ede4_u0<=reg_7a0a4746_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_34313572_u0<=1'h0;
else reg_34313572_u0<=reg_319759b9_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_328d47c8_u0<=1'h0;
else reg_328d47c8_u0<=reg_6ee42c26_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3bf5fabd_u0<=1'h0;
else reg_3bf5fabd_u0<=reg_5df5aff9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_27394bed_result_delayed_u0<=1'h0;
else reg_27394bed_result_delayed_u0<=reg_27394bed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_107de137_u0<=1'h0;
else reg_107de137_u0<=reg_0dcebdfe_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a0a4746_u0<=1'h0;
else reg_7a0a4746_u0<=reg_73231fe1_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_561bf6ff_result_delayed_u0<=1'h0;
else reg_561bf6ff_result_delayed_u0<=reg_561bf6ff_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_58245975_u0<=1'h0;
else reg_58245975_u0<=reg_723816cc_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2913cc47_u0<=1'h0;
else reg_2913cc47_u0<=reg_49eb7136_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_41757d04_result_delayed_result_delayed_u0<=1'h0;
else reg_41757d04_result_delayed_result_delayed_u0<=reg_41757d04_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_27cdb75f_result_delayed_u0<=1'h0;
else reg_27cdb75f_result_delayed_u0<=reg_27cdb75f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_107de137_result_delayed_u0<=1'h0;
else reg_107de137_result_delayed_u0<=reg_107de137_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0ffd27c0_result_delayed_u0<=1'h0;
else reg_0ffd27c0_result_delayed_u0<=reg_0ffd27c0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_44a091fd_u0<=1'h0;
else reg_44a091fd_u0<=reg_4b2b9289_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_30bea5e3_u0<=1'h0;
else reg_30bea5e3_u0<=reg_0178db0e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2fe8a6b5_u0<=1'h0;
else reg_2fe8a6b5_u0<=reg_4692efed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_55d7a1ff_result_delayed_result_delayed_u0<=1'h0;
else reg_55d7a1ff_result_delayed_result_delayed_u0<=reg_55d7a1ff_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3ac9d797_u0<=1'h0;
else reg_3ac9d797_u0<=reg_619a949e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_635d5720_result_delayed_u0<=1'h0;
else reg_635d5720_result_delayed_u0<=reg_635d5720_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2913cc47_result_delayed_u0<=1'h0;
else reg_2913cc47_result_delayed_u0<=reg_2913cc47_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_306c2418_result_delayed_u0<=1'h0;
else reg_306c2418_result_delayed_u0<=reg_306c2418_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4e506b37_u0<=1'h0;
else reg_4e506b37_u0<=reg_4cd5885f_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_27faaa92_u0<=1'h0;
else reg_27faaa92_u0<=reg_3bf5fabd_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_107de137_result_delayed_result_delayed_u0<=1'h0;
else reg_107de137_result_delayed_result_delayed_u0<=reg_107de137_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_31f84093_u0<=1'h0;
else reg_31f84093_u0<=reg_561ae0f2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_247a1111_u0<=1'h0;
else reg_247a1111_u0<=reg_5d3a8c49_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2fe8a6b5_result_delayed_u0<=1'h0;
else reg_2fe8a6b5_result_delayed_u0<=reg_2fe8a6b5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4a382354_u0<=1'h0;
else reg_4a382354_u0<=reg_0c928251_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6b0d2e60_u0<=1'h0;
else reg_6b0d2e60_u0<=reg_343bd27c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5cbbf0a1_result_delayed_u0<=1'h0;
else reg_5cbbf0a1_result_delayed_u0<=reg_5cbbf0a1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a0a4746_result_delayed_u0<=1'h0;
else reg_7a0a4746_result_delayed_u0<=reg_7a0a4746_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_619a949e_result_delayed_u0<=1'h0;
else reg_619a949e_result_delayed_u0<=reg_619a949e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5d3a8c49_u0<=1'h0;
else reg_5d3a8c49_u0<=reg_1eb746e3_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3d110516_result_delayed_u0<=1'h0;
else reg_3d110516_result_delayed_u0<=reg_3d110516_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_35c048b4_u0<=1'h0;
else reg_35c048b4_u0<=reg_7368e3a4_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_49eb7136_result_delayed_u0<=1'h0;
else reg_49eb7136_result_delayed_u0<=reg_49eb7136_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_213ddd8e_result_delayed_u0<=1'h0;
else reg_213ddd8e_result_delayed_u0<=reg_213ddd8e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7c5e9123_u0<=1'h0;
else reg_7c5e9123_u0<=reg_27394bed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4692efed_u0<=1'h0;
else reg_4692efed_u0<=reg_4bda7e7a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_166d6bed_u0<=1'h0;
else reg_166d6bed_u0<=reg_63d04af9_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_47d1d653_u0<=1'h0;
else reg_47d1d653_u0<=reg_7984ac77_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_13e88a6a_u0<=1'h0;
else reg_13e88a6a_u0<=reg_7bb0f302_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_79dd91a5_result_delayed_u0<=1'h0;
else reg_79dd91a5_result_delayed_u0<=reg_79dd91a5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_14ebcd6f_u0<=1'h0;
else reg_14ebcd6f_u0<=reg_2159053d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_157eb4fb_u0<=1'h0;
else reg_157eb4fb_u0<=reg_0ba46dcc_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_32992b13_u0<=1'h0;
else reg_32992b13_u0<=reg_00c68dc2_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1e3be3b6_u0<=1'h0;
else reg_1e3be3b6_u0<=reg_3771f97a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7ec5534b_u0<=1'h0;
else reg_7ec5534b_u0<=reg_0da90157_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0d8e6001_u0<=1'h0;
else reg_0d8e6001_u0<=reg_31278190_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4cd5885f_result_delayed_result_delayed_u0<=1'h0;
else reg_4cd5885f_result_delayed_result_delayed_u0<=reg_4cd5885f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_03bb9a29_u0<=1'h0;
else reg_03bb9a29_u0<=reg_4cdea096_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_50412dd3_u0<=1'h0;
else reg_50412dd3_u0<=reg_4bf77a1c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_322587b0_u0<=1'h0;
else reg_322587b0_u0<=reg_7432549f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3a122388_u0<=1'h0;
else reg_3a122388_u0<=reg_7b860f51_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1f4a72d1_u0<=1'h0;
else reg_1f4a72d1_u0<=reg_65390362_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_398e1010_u0<=1'h0;
else reg_398e1010_u0<=reg_1d5ae331_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4bda7e7a_u0<=1'h0;
else reg_4bda7e7a_u0<=reg_50e04075_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6b0d2e60_result_delayed_u0<=1'h0;
else reg_6b0d2e60_result_delayed_u0<=reg_6b0d2e60_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4b2b9289_u0<=1'h0;
else reg_4b2b9289_u0<=reg_3cd29fd9_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_40236581_u0<=1'h0;
else reg_40236581_u0<=reg_01f9b917_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7203dba7_u0<=1'h0;
else reg_7203dba7_u0<=reg_37c4aa7f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_507b6cf9_result_delayed_u0<=1'h0;
else reg_507b6cf9_result_delayed_u0<=reg_507b6cf9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6e4f17e9_u0<=1'h0;
else reg_6e4f17e9_u0<=reg_414b944f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_12e5bf43_u0<=1'h0;
else reg_12e5bf43_u0<=reg_5367bbad_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4f83ce24_u0<=1'h0;
else reg_4f83ce24_u0<=reg_608e408d_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_774d2b58_result_delayed_u0<=1'h0;
else reg_774d2b58_result_delayed_u0<=reg_774d2b58_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01f9b917_result_delayed_u0<=1'h0;
else reg_01f9b917_result_delayed_u0<=reg_01f9b917_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_776a1f94_result_delayed_u0<=1'h0;
else reg_776a1f94_result_delayed_u0<=reg_776a1f94_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_490168aa_u0<=1'h0;
else reg_490168aa_u0<=reg_103f4835_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4bda7e7a_result_delayed_u0<=1'h0;
else reg_4bda7e7a_result_delayed_u0<=reg_4bda7e7a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5c0a547e_result_delayed_result_delayed_u0<=1'h0;
else reg_5c0a547e_result_delayed_result_delayed_u0<=reg_5c0a547e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6cdc1173_u0<=1'h0;
else reg_6cdc1173_u0<=reg_36d51882_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5367bbad_result_delayed_u0<=1'h0;
else reg_5367bbad_result_delayed_u0<=reg_5367bbad_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3365b2d6_u0<=1'h0;
else reg_3365b2d6_u0<=reg_5cbbf0a1_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_78922926_u0<=1'h0;
else reg_78922926_u0<=reg_2b4cee92_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4a747bcd_u0<=1'h0;
else reg_4a747bcd_u0<=reg_02179ae1_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_37c4aa7f_u0<=1'h0;
else reg_37c4aa7f_u0<=reg_156fe33d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_73231fe1_result_delayed_u0<=1'h0;
else reg_73231fe1_result_delayed_u0<=reg_73231fe1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_33bcd31f_result_delayed_u0<=1'h0;
else reg_33bcd31f_result_delayed_u0<=reg_33bcd31f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1ba8b669_u0<=1'h0;
else reg_1ba8b669_u0<=reg_08701441_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4fd02acb_result_delayed_u0<=1'h0;
else reg_4fd02acb_result_delayed_u0<=reg_4fd02acb_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_35bbb476_u0<=1'h0;
else reg_35bbb476_u0<=reg_6f9f0292_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_720d5fdc_u0<=1'h0;
else reg_720d5fdc_u0<=reg_3d3b97a5_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0f95e647_u0<=1'h0;
else reg_0f95e647_u0<=reg_56d52bdd_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5d1c80c9_u0<=1'h0;
else reg_5d1c80c9_u0<=reg_559271a8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_63d04af9_result_delayed_u0<=1'h0;
else reg_63d04af9_result_delayed_u0<=reg_63d04af9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2b4cee92_u0<=1'h0;
else reg_2b4cee92_u0<=reg_1afd62a7_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_20599c2d_result_delayed_u0<=1'h0;
else reg_20599c2d_result_delayed_u0<=reg_20599c2d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5c6cbd8d_u0<=1'h0;
else reg_5c6cbd8d_u0<=reg_7c5e9123_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_07979748_result_delayed_u0<=1'h0;
else reg_07979748_result_delayed_u0<=reg_07979748_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7368e3a4_result_delayed_u0<=1'h0;
else reg_7368e3a4_result_delayed_u0<=reg_7368e3a4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1fa5dbf4_result_delayed_u0<=1'h0;
else reg_1fa5dbf4_result_delayed_u0<=reg_1fa5dbf4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1bd6ae3f_u0<=1'h0;
else reg_1bd6ae3f_u0<=reg_5eb4b0ba_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4bf77a1c_u0<=1'h0;
else reg_4bf77a1c_u0<=reg_2fe8a6b5_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_771e534d_result_delayed_u0<=1'h0;
else reg_771e534d_result_delayed_u0<=reg_771e534d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_25c1902c_u0<=1'h0;
else reg_25c1902c_u0<=reg_1e3be3b6_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_68fe950f_u0<=1'h0;
else reg_68fe950f_u0<=reg_64544e65_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7984ac77_u0<=1'h0;
else reg_7984ac77_u0<=reg_796d6b70_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_32797234_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_32797234_result_delayed_result_delayed_result_delayed_u0<=reg_32797234_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7b860f51_result_delayed_u0<=1'h0;
else reg_7b860f51_result_delayed_u0<=reg_7b860f51_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_58245975_result_delayed_u0<=1'h0;
else reg_58245975_result_delayed_u0<=reg_58245975_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_626c9aa9_result_delayed_u0<=1'h0;
else reg_626c9aa9_result_delayed_u0<=reg_626c9aa9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_728582a2_result_delayed_u0<=1'h0;
else reg_728582a2_result_delayed_u0<=reg_728582a2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_04257c62_result_delayed_u0<=1'h0;
else reg_04257c62_result_delayed_u0<=reg_04257c62_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4262839e_u0<=1'h0;
else reg_4262839e_u0<=reg_43d7d4e5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_74845d78_u0<=1'h0;
else reg_74845d78_u0<=reg_3601783e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_248ca170_u0<=1'h0;
else reg_248ca170_u0<=reg_03167f2b_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0dcebdfe_result_delayed_u0<=1'h0;
else reg_0dcebdfe_result_delayed_u0<=reg_0dcebdfe_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_41757d04_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_41757d04_result_delayed_result_delayed_result_delayed_u0<=reg_41757d04_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2e9b949b_u0<=1'h0;
else reg_2e9b949b_u0<=reg_247a1111_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_739d919c_u0<=1'h0;
else reg_739d919c_u0<=reg_78922926_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_12e5bf43_result_delayed_u0<=1'h0;
else reg_12e5bf43_result_delayed_u0<=reg_12e5bf43_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0629ba72_result_delayed_u0<=1'h0;
else reg_0629ba72_result_delayed_u0<=reg_0629ba72_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6da911c6_result_delayed_u0<=1'h0;
else reg_6da911c6_result_delayed_u0<=reg_6da911c6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_43dfbb10_result_delayed_u0<=1'h0;
else reg_43dfbb10_result_delayed_u0<=reg_43dfbb10_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_776a1f94_result_delayed_result_delayed_u0<=1'h0;
else reg_776a1f94_result_delayed_result_delayed_u0<=reg_776a1f94_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a0a4746_result_delayed_result_delayed_u0<=1'h0;
else reg_7a0a4746_result_delayed_result_delayed_u0<=reg_7a0a4746_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3771f97a_u0<=1'h0;
else reg_3771f97a_u0<=reg_6da911c6_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_248ca170_result_delayed_u0<=1'h0;
else reg_248ca170_result_delayed_u0<=reg_248ca170_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5df5aff9_u0<=1'h0;
else reg_5df5aff9_u0<=reg_0e249eb7_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5eb4b0ba_u0<=1'h0;
else reg_5eb4b0ba_u0<=reg_25c1902c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2b82898d_u0<=1'h0;
else reg_2b82898d_u0<=reg_248ca170_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4692efed_result_delayed_u0<=1'h0;
else reg_4692efed_result_delayed_u0<=reg_4692efed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_559271a8_result_delayed_u0<=1'h0;
else reg_559271a8_result_delayed_u0<=reg_559271a8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_723816cc_result_delayed_u0<=1'h0;
else reg_723816cc_result_delayed_u0<=reg_723816cc_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_05d67bc0_u0<=1'h0;
else reg_05d67bc0_u0<=reg_74845d78_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6ee280fb_u0<=1'h0;
else reg_6ee280fb_u0<=reg_3c50f618_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a591648_result_delayed_u0<=1'h0;
else reg_7a591648_result_delayed_u0<=reg_7a591648_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_796d6b70_u0<=1'h0;
else reg_796d6b70_u0<=reg_10ae20df_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6da911c6_result_delayed_result_delayed_u0<=1'h0;
else reg_6da911c6_result_delayed_result_delayed_u0<=reg_6da911c6_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3562c342_u0<=1'h0;
else reg_3562c342_u0<=reg_43dfbb10_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5cbbf0a1_result_delayed_result_delayed_u0<=1'h0;
else reg_5cbbf0a1_result_delayed_result_delayed_u0<=reg_5cbbf0a1_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_35875fa3_u0<=1'h0;
else reg_35875fa3_u0<=reg_07979748_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_328d47c8_result_delayed_u0<=1'h0;
else reg_328d47c8_result_delayed_u0<=reg_328d47c8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4cdea096_result_delayed_u0<=1'h0;
else reg_4cdea096_result_delayed_u0<=reg_4cdea096_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_103f4835_result_delayed_u0<=1'h0;
else reg_103f4835_result_delayed_u0<=reg_103f4835_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1204a325_result_delayed_u0<=1'h0;
else reg_1204a325_result_delayed_u0<=reg_1204a325_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_64544e65_u0<=1'h0;
else reg_64544e65_u0<=reg_655155f8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_655155f8_result_delayed_u0<=1'h0;
else reg_655155f8_result_delayed_u0<=reg_655155f8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_31278190_result_delayed_u0<=1'h0;
else reg_31278190_result_delayed_u0<=reg_31278190_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_27410d75_u0<=1'h0;
else reg_27410d75_u0<=and_u1764_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_579fa5aa_u0<=1'h0;
else reg_579fa5aa_u0<=reg_4262839e_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1e3be3b6_result_delayed_u0<=1'h0;
else reg_1e3be3b6_result_delayed_u0<=reg_1e3be3b6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_02d9964d_result_delayed_u0<=1'h0;
else reg_02d9964d_result_delayed_u0<=reg_02d9964d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4db5d9f8_result_delayed_u0<=1'h0;
else reg_4db5d9f8_result_delayed_u0<=reg_4db5d9f8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3601783e_u0<=1'h0;
else reg_3601783e_u0<=reg_42f3b02c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_08701441_result_delayed_u0<=1'h0;
else reg_08701441_result_delayed_u0<=reg_08701441_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_066f602e_u0<=1'h0;
else reg_066f602e_u0<=reg_3dfa0f2c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_19f2d151_result_delayed_u0<=1'h0;
else reg_19f2d151_result_delayed_u0<=reg_19f2d151_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7c98e992_result_delayed_u0<=1'h0;
else reg_7c98e992_result_delayed_u0<=reg_7c98e992_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7c9a16d9_u0<=1'h0;
else reg_7c9a16d9_u0<=reg_02d9964d_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_343bd27c_u0<=1'h0;
else reg_343bd27c_u0<=reg_561bf6ff_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2b1f6158_u0<=1'h0;
else reg_2b1f6158_u0<=reg_6e4f17e9_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3c50f618_u0<=1'h0;
else reg_3c50f618_u0<=reg_5e49be57_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3bf5fabd_result_delayed_u0<=1'h0;
else reg_3bf5fabd_result_delayed_u0<=reg_3bf5fabd_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7c5e9123_result_delayed_u0<=1'h0;
else reg_7c5e9123_result_delayed_u0<=reg_7c5e9123_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_156fe33d_u0<=1'h0;
else reg_156fe33d_u0<=reg_2c6d2fd0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4cdea096_result_delayed_result_delayed_u0<=1'h0;
else reg_4cdea096_result_delayed_result_delayed_u0<=reg_4cdea096_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_14ebcd6f_result_delayed_u0<=1'h0;
else reg_14ebcd6f_result_delayed_u0<=reg_14ebcd6f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_170037b2_result_delayed_u0<=1'h0;
else reg_170037b2_result_delayed_u0<=reg_170037b2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_30e53c09_result_delayed_u0<=1'h0;
else reg_30e53c09_result_delayed_u0<=reg_30e53c09_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6fa9d1fe_u0<=1'h0;
else reg_6fa9d1fe_u0<=reg_0ef60446_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_36d51882_u0<=1'h0;
else reg_36d51882_u0<=reg_6d11391e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4262839e_result_delayed_u0<=1'h0;
else reg_4262839e_result_delayed_u0<=reg_4262839e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_65390362_u0<=1'h0;
else reg_65390362_u0<=reg_0da887c4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00c68dc2_result_delayed_u0<=1'h0;
else reg_00c68dc2_result_delayed_u0<=reg_00c68dc2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6f9f0292_result_delayed_u0<=1'h0;
else reg_6f9f0292_result_delayed_u0<=reg_6f9f0292_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2711b972_u0<=1'h0;
else reg_2711b972_u0<=reg_2eee6ac6_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_33bcd31f_result_delayed_result_delayed_u0<=1'h0;
else reg_33bcd31f_result_delayed_result_delayed_u0<=reg_33bcd31f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2eee6ac6_result_delayed_result_delayed_u0<=1'h0;
else reg_2eee6ac6_result_delayed_result_delayed_u0<=reg_2eee6ac6_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_357d771a_u0<=1'h0;
else reg_357d771a_u0<=reg_7080240a_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5bf74d9f_u0<=1'h0;
else reg_5bf74d9f_u0<=reg_71343346_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0ba46dcc_u0<=1'h0;
else reg_0ba46dcc_u0<=reg_6bb9ab9e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7d792c42_result_delayed_u0<=1'h0;
else reg_7d792c42_result_delayed_u0<=reg_7d792c42_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_772bbfa5_result_delayed_u0<=1'h0;
else reg_772bbfa5_result_delayed_u0<=reg_772bbfa5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1d5ae331_u0<=1'h0;
else reg_1d5ae331_u0<=reg_73b33bd3_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0da887c4_u0<=1'h0;
else reg_0da887c4_u0<=reg_23b89b62_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_32301a2a_result_delayed_result_delayed_u0<=1'h0;
else reg_32301a2a_result_delayed_result_delayed_u0<=reg_32301a2a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_41a8efc6_u0<=1'h0;
else reg_41a8efc6_u0<=reg_69761137_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7bb0f302_result_delayed_u0<=1'h0;
else reg_7bb0f302_result_delayed_u0<=reg_7bb0f302_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6bb9ab9e_result_delayed_u0<=1'h0;
else reg_6bb9ab9e_result_delayed_u0<=reg_6bb9ab9e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_71343346_u0<=1'h0;
else reg_71343346_u0<=reg_2586ddf0_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2f9c95e8_u0<=1'h0;
else reg_2f9c95e8_u0<=reg_7a591648_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0178db0e_u0<=1'h0;
else reg_0178db0e_u0<=reg_5c0a547e_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5eb4b0ba_result_delayed_u0<=1'h0;
else reg_5eb4b0ba_result_delayed_u0<=reg_5eb4b0ba_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_02d9964d_result_delayed_result_delayed_u0<=1'h0;
else reg_02d9964d_result_delayed_result_delayed_u0<=reg_02d9964d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_27394bed_result_delayed_result_delayed_u0<=1'h0;
else reg_27394bed_result_delayed_result_delayed_u0<=reg_27394bed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_68fe950f_result_delayed_u0<=1'h0;
else reg_68fe950f_result_delayed_u0<=reg_68fe950f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7bb0f302_result_delayed_result_delayed_u0<=1'h0;
else reg_7bb0f302_result_delayed_result_delayed_u0<=reg_7bb0f302_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_45429118_result_delayed_u0<=1'h0;
else reg_45429118_result_delayed_u0<=reg_45429118_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_19f2d151_result_delayed_result_delayed_u0<=1'h0;
else reg_19f2d151_result_delayed_result_delayed_u0<=reg_19f2d151_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_32992b13_result_delayed_u0<=1'h0;
else reg_32992b13_result_delayed_u0<=reg_32992b13_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_10ae20df_result_delayed_result_delayed_u0<=1'h0;
else reg_10ae20df_result_delayed_result_delayed_u0<=reg_10ae20df_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1e3be3b6_result_delayed_result_delayed_u0<=1'h0;
else reg_1e3be3b6_result_delayed_result_delayed_u0<=reg_1e3be3b6_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_56d52bdd_result_delayed_u0<=1'h0;
else reg_56d52bdd_result_delayed_u0<=reg_56d52bdd_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6b0d2e60_result_delayed_result_delayed_u0<=1'h0;
else reg_6b0d2e60_result_delayed_result_delayed_u0<=reg_6b0d2e60_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a230a1a_result_delayed_u0<=1'h0;
else reg_7a230a1a_result_delayed_u0<=reg_7a230a1a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0ba46dcc_result_delayed_u0<=1'h0;
else reg_0ba46dcc_result_delayed_u0<=reg_0ba46dcc_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_247e36e9_u0<=1'h0;
else reg_247e36e9_u0<=reg_31f84093_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_248ca170_result_delayed_result_delayed_u0<=1'h0;
else reg_248ca170_result_delayed_result_delayed_u0<=reg_248ca170_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_43dfbb10_result_delayed_result_delayed_u0<=1'h0;
else reg_43dfbb10_result_delayed_result_delayed_u0<=reg_43dfbb10_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_490168aa_result_delayed_u0<=1'h0;
else reg_490168aa_result_delayed_u0<=reg_490168aa_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4cd5885f_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_4cd5885f_result_delayed_result_delayed_result_delayed_u0<=reg_4cd5885f_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4262839e_result_delayed_result_delayed_u0<=1'h0;
else reg_4262839e_result_delayed_result_delayed_u0<=reg_4262839e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_31f84093_result_delayed_u0<=1'h0;
else reg_31f84093_result_delayed_u0<=reg_31f84093_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3d3b97a5_u0<=1'h0;
else reg_3d3b97a5_u0<=reg_157eb4fb_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_02179ae1_result_delayed_u0<=1'h0;
else reg_02179ae1_result_delayed_u0<=reg_02179ae1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_561bf6ff_result_delayed_result_delayed_u0<=1'h0;
else reg_561bf6ff_result_delayed_result_delayed_u0<=reg_561bf6ff_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_03167f2b_result_delayed_result_delayed_u0<=1'h0;
else reg_03167f2b_result_delayed_result_delayed_u0<=reg_03167f2b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4ce52437_result_delayed_u0<=1'h0;
else reg_4ce52437_result_delayed_u0<=reg_4ce52437_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_19f2d151_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_19f2d151_result_delayed_result_delayed_result_delayed_u0<=reg_19f2d151_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6ca7ede4_result_delayed_u0<=1'h0;
else reg_6ca7ede4_result_delayed_u0<=reg_6ca7ede4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0ef60446_u0<=1'h0;
else reg_0ef60446_u0<=reg_297e0532_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2fe8a6b5_result_delayed_result_delayed_u0<=1'h0;
else reg_2fe8a6b5_result_delayed_result_delayed_u0<=reg_2fe8a6b5_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6ff27b40_result_delayed_u0<=1'h0;
else reg_6ff27b40_result_delayed_u0<=reg_6ff27b40_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4cdea096_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_4cdea096_result_delayed_result_delayed_result_delayed_u0<=reg_4cdea096_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5cbbf0a1_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_5cbbf0a1_result_delayed_result_delayed_result_delayed_u0<=reg_5cbbf0a1_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7432549f_result_delayed_u0<=1'h0;
else reg_7432549f_result_delayed_u0<=reg_7432549f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6ee42c26_u0<=1'h0;
else reg_6ee42c26_u0<=reg_776a1f94_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4692efed_result_delayed_result_delayed_u0<=1'h0;
else reg_4692efed_result_delayed_result_delayed_u0<=reg_4692efed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0c928251_u0<=1'h0;
else reg_0c928251_u0<=reg_22387d0e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_20599c2d_result_delayed_result_delayed_u0<=1'h0;
else reg_20599c2d_result_delayed_result_delayed_u0<=reg_20599c2d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_319759b9_result_delayed_u0<=1'h0;
else reg_319759b9_result_delayed_u0<=reg_319759b9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_62251200_result_delayed_u0<=1'h0;
else reg_62251200_result_delayed_u0<=reg_62251200_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7d792c42_result_delayed_result_delayed_u0<=1'h0;
else reg_7d792c42_result_delayed_result_delayed_u0<=reg_7d792c42_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1fa5dbf4_result_delayed_result_delayed_u0<=1'h0;
else reg_1fa5dbf4_result_delayed_result_delayed_u0<=reg_1fa5dbf4_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5eb4b0ba_result_delayed_result_delayed_u0<=1'h0;
else reg_5eb4b0ba_result_delayed_result_delayed_u0<=reg_5eb4b0ba_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3dfa0f2c_u0<=1'h0;
else reg_3dfa0f2c_u0<=reg_22e2922b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_55d7a1ff_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_55d7a1ff_result_delayed_result_delayed_result_delayed_u0<=reg_55d7a1ff_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6ee42c26_result_delayed_u0<=1'h0;
else reg_6ee42c26_result_delayed_u0<=reg_6ee42c26_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_26bc9067_u0<=1'h0;
else reg_26bc9067_u0<=reg_3d110516_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1ba8b669_result_delayed_u0<=1'h0;
else reg_1ba8b669_result_delayed_u0<=reg_1ba8b669_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3d75c9ae_result_delayed_u0<=1'h0;
else reg_3d75c9ae_result_delayed_u0<=reg_3d75c9ae_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_31f84093_result_delayed_result_delayed_u0<=1'h0;
else reg_31f84093_result_delayed_result_delayed_u0<=reg_31f84093_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_42f3b02c_u0<=1'h0;
else reg_42f3b02c_u0<=reg_326d6def_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2afa8c1b_u0<=1'h0;
else reg_2afa8c1b_u0<=reg_579fa5aa_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7c5e9123_result_delayed_result_delayed_u0<=1'h0;
else reg_7c5e9123_result_delayed_result_delayed_u0<=reg_7c5e9123_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2ab2a055_u0<=1'h0;
else reg_2ab2a055_u0<=and_u1765_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_69761137_result_delayed_u0<=1'h0;
else reg_69761137_result_delayed_u0<=reg_69761137_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_561ae0f2_u0<=1'h0;
else reg_561ae0f2_u0<=reg_44cb88e0_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1eb746e3_result_delayed_u0<=1'h0;
else reg_1eb746e3_result_delayed_u0<=reg_1eb746e3_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_10ff65be_result_delayed_u0<=1'h0;
else reg_10ff65be_result_delayed_u0<=reg_10ff65be_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4e506b37_result_delayed_u0<=1'h0;
else reg_4e506b37_result_delayed_u0<=reg_4e506b37_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3a122388_result_delayed_u0<=1'h0;
else reg_3a122388_result_delayed_u0<=reg_3a122388_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_31f84093_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_31f84093_result_delayed_result_delayed_result_delayed_u0<=reg_31f84093_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0ae85810_u0<=1'h0;
else reg_0ae85810_u0<=reg_40236581_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3c50f618_result_delayed_u0<=1'h0;
else reg_3c50f618_result_delayed_u0<=reg_3c50f618_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4692efed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_4692efed_result_delayed_result_delayed_result_delayed_u0<=reg_4692efed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6f6443d2_result_delayed_u0<=1'h0;
else reg_6f6443d2_result_delayed_u0<=reg_6f6443d2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4d69442a_result_delayed_u0<=1'h0;
else reg_4d69442a_result_delayed_u0<=reg_4d69442a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3cd29fd9_u0<=1'h0;
else reg_3cd29fd9_u0<=reg_3ac9d797_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_73b33bd3_result_delayed_u0<=1'h0;
else reg_73b33bd3_result_delayed_u0<=reg_73b33bd3_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_25c1902c_result_delayed_u0<=1'h0;
else reg_25c1902c_result_delayed_u0<=reg_25c1902c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_729e0d87_u0<=1'h0;
else reg_729e0d87_u0<=reg_72f7e7fe_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_30bea5e3_result_delayed_u0<=1'h0;
else reg_30bea5e3_result_delayed_u0<=reg_30bea5e3_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_44cb88e0_result_delayed_u0<=1'h0;
else reg_44cb88e0_result_delayed_u0<=reg_44cb88e0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_606de772_u0<=1'h0;
else reg_606de772_u0<=reg_4bc0004f_result_delayed_u0;
end
assign and_u1764_u0=and_u1760_u0&and_u1767_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_71343346_result_delayed_u0<=1'h0;
else reg_71343346_result_delayed_u0<=reg_71343346_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_49eb7136_result_delayed_result_delayed_u0<=1'h0;
else reg_49eb7136_result_delayed_result_delayed_u0<=reg_49eb7136_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2586ddf0_result_delayed_result_delayed_u0<=1'h0;
else reg_2586ddf0_result_delayed_result_delayed_u0<=reg_2586ddf0_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7352b877_u0<=1'h0;
else reg_7352b877_u0<=reg_09fdcdde_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_40236581_result_delayed_u0<=1'h0;
else reg_40236581_result_delayed_u0<=reg_40236581_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_414b944f_result_delayed_u0<=1'h0;
else reg_414b944f_result_delayed_u0<=reg_414b944f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_739d919c_result_delayed_u0<=1'h0;
else reg_739d919c_result_delayed_u0<=reg_739d919c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3cd29fd9_result_delayed_u0<=1'h0;
else reg_3cd29fd9_result_delayed_u0<=reg_3cd29fd9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_188534c8_result_delayed_u0<=1'h0;
else reg_188534c8_result_delayed_u0<=reg_188534c8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_09fdcdde_result_delayed_u0<=1'h0;
else reg_09fdcdde_result_delayed_u0<=reg_09fdcdde_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_43d7d4e5_u0<=1'h0;
else reg_43d7d4e5_u0<=reg_1e307217_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_02179ae1_result_delayed_result_delayed_u0<=1'h0;
else reg_02179ae1_result_delayed_result_delayed_u0<=reg_02179ae1_result_delayed_u0;
end
assign mux_u180=(and_u1765_u0)?1'h1:1'h0;
assign or_u482_u0=and_u1765_u0|and_u1763_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_22387d0e_u0<=1'h0;
else reg_22387d0e_u0<=reg_635d5720_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_32301a2a_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_32301a2a_result_delayed_result_delayed_result_delayed_u0<=reg_32301a2a_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_357d771a_result_delayed_u0<=1'h0;
else reg_357d771a_result_delayed_u0<=reg_357d771a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5e49be57_result_delayed_u0<=1'h0;
else reg_5e49be57_result_delayed_u0<=reg_5e49be57_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_776a1f94_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_776a1f94_result_delayed_result_delayed_result_delayed_u0<=reg_776a1f94_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_552e2e6e_u0<=1'h0;
else reg_552e2e6e_u0<=reg_4e506b37_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2711b972_result_delayed_u0<=1'h0;
else reg_2711b972_result_delayed_u0<=reg_2711b972_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_398e1010_result_delayed_u0<=1'h0;
else reg_398e1010_result_delayed_u0<=reg_398e1010_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_78922926_result_delayed_u0<=1'h0;
else reg_78922926_result_delayed_u0<=reg_78922926_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_630a4c43_u0<=1'h0;
else reg_630a4c43_u0<=reg_16db469f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4939b9f8_result_delayed_u0<=1'h0;
else reg_4939b9f8_result_delayed_u0<=reg_4939b9f8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0da90157_result_delayed_u0<=1'h0;
else reg_0da90157_result_delayed_u0<=reg_0da90157_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_635d5720_result_delayed_result_delayed_u0<=1'h0;
else reg_635d5720_result_delayed_result_delayed_u0<=reg_635d5720_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_343bd27c_result_delayed_u0<=1'h0;
else reg_343bd27c_result_delayed_u0<=reg_343bd27c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3e0fda11_result_delayed_u0<=1'h0;
else reg_3e0fda11_result_delayed_u0<=reg_3e0fda11_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3ac9d797_result_delayed_u0<=1'h0;
else reg_3ac9d797_result_delayed_u0<=reg_3ac9d797_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3d3b97a5_result_delayed_u0<=1'h0;
else reg_3d3b97a5_result_delayed_u0<=reg_3d3b97a5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3562c342_result_delayed_u0<=1'h0;
else reg_3562c342_result_delayed_u0<=reg_3562c342_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_157eb4fb_result_delayed_u0<=1'h0;
else reg_157eb4fb_result_delayed_u0<=reg_157eb4fb_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6ccfd5e8_result_delayed_u0<=1'h0;
else reg_6ccfd5e8_result_delayed_u0<=reg_6ccfd5e8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2b2ea879_u0<=1'h0;
else reg_2b2ea879_u0<=reg_55d7a1ff_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_02179ae1_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_02179ae1_result_delayed_result_delayed_result_delayed_u0<=reg_02179ae1_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_626c9aa9_result_delayed_result_delayed_u0<=1'h0;
else reg_626c9aa9_result_delayed_result_delayed_u0<=reg_626c9aa9_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4e506b37_result_delayed_result_delayed_u0<=1'h0;
else reg_4e506b37_result_delayed_result_delayed_u0<=reg_4e506b37_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2159053d_result_delayed_u0<=1'h0;
else reg_2159053d_result_delayed_u0<=reg_2159053d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7ec5534b_result_delayed_u0<=1'h0;
else reg_7ec5534b_result_delayed_u0<=reg_7ec5534b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0ffd27c0_result_delayed_result_delayed_u0<=1'h0;
else reg_0ffd27c0_result_delayed_result_delayed_u0<=reg_0ffd27c0_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_32797234_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_32797234_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_32797234_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3d110516_result_delayed_result_delayed_u0<=1'h0;
else reg_3d110516_result_delayed_result_delayed_u0<=reg_3d110516_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7080240a_result_delayed_result_delayed_u0<=1'h0;
else reg_7080240a_result_delayed_result_delayed_u0<=reg_7080240a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_55d7a1ff_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_55d7a1ff_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_55d7a1ff_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6ca7ede4_result_delayed_result_delayed_u0<=1'h0;
else reg_6ca7ede4_result_delayed_result_delayed_u0<=reg_6ca7ede4_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_23b89b62_result_delayed_u0<=1'h0;
else reg_23b89b62_result_delayed_u0<=reg_23b89b62_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1afd62a7_result_delayed_u0<=1'h0;
else reg_1afd62a7_result_delayed_u0<=reg_1afd62a7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_35875fa3_result_delayed_u0<=1'h0;
else reg_35875fa3_result_delayed_u0<=reg_35875fa3_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_579fa5aa_result_delayed_u0<=1'h0;
else reg_579fa5aa_result_delayed_u0<=reg_579fa5aa_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2e3a4ef5_result_delayed_result_delayed_u0<=1'h0;
else reg_2e3a4ef5_result_delayed_result_delayed_u0<=reg_2e3a4ef5_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_772bbfa5_result_delayed_result_delayed_u0<=1'h0;
else reg_772bbfa5_result_delayed_result_delayed_u0<=reg_772bbfa5_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_50e04075_result_delayed_u0<=1'h0;
else reg_50e04075_result_delayed_u0<=reg_50e04075_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1bd6ae3f_result_delayed_u0<=1'h0;
else reg_1bd6ae3f_result_delayed_u0<=reg_1bd6ae3f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_326d6def_u0<=1'h0;
else reg_326d6def_u0<=reg_6ee280fb_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6e4f17e9_result_delayed_u0<=1'h0;
else reg_6e4f17e9_result_delayed_u0<=reg_6e4f17e9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_608e408d_result_delayed_result_delayed_u0<=1'h0;
else reg_608e408d_result_delayed_result_delayed_u0<=reg_608e408d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7d792c42_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_7d792c42_result_delayed_result_delayed_result_delayed_u0<=reg_7d792c42_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_066f602e_result_delayed_u0<=1'h0;
else reg_066f602e_result_delayed_u0<=reg_066f602e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2a9c2111_u0<=1'h0;
else reg_2a9c2111_u0<=reg_3a122388_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_248ca170_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_248ca170_result_delayed_result_delayed_result_delayed_u0<=reg_248ca170_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6da911c6_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_6da911c6_result_delayed_result_delayed_result_delayed_u0<=reg_6da911c6_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4bc0004f_u0<=1'h0;
else reg_4bc0004f_u0<=reg_04257c62_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_04257c62_result_delayed_result_delayed_u0<=1'h0;
else reg_04257c62_result_delayed_result_delayed_u0<=reg_04257c62_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3a122388_result_delayed_result_delayed_u0<=1'h0;
else reg_3a122388_result_delayed_result_delayed_u0<=reg_3a122388_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_056e42f2_u0<=1'h0;
else reg_056e42f2_u0<=reg_30bea5e3_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_319759b9_result_delayed_result_delayed_u0<=1'h0;
else reg_319759b9_result_delayed_result_delayed_u0<=reg_319759b9_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4db5d9f8_result_delayed_result_delayed_u0<=1'h0;
else reg_4db5d9f8_result_delayed_result_delayed_u0<=reg_4db5d9f8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_510951b8_result_delayed_u0<=1'h0;
else reg_510951b8_result_delayed_u0<=reg_510951b8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_22e2922b_result_delayed_u0<=1'h0;
else reg_22e2922b_result_delayed_u0<=reg_22e2922b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6d11391e_result_delayed_u0<=1'h0;
else reg_6d11391e_result_delayed_u0<=reg_6d11391e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1e307217_result_delayed_u0<=1'h0;
else reg_1e307217_result_delayed_u0<=reg_1e307217_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2b82898d_result_delayed_u0<=1'h0;
else reg_2b82898d_result_delayed_u0<=reg_2b82898d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1d5ae331_result_delayed_u0<=1'h0;
else reg_1d5ae331_result_delayed_u0<=reg_1d5ae331_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_41757d04_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_41757d04_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_41757d04_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_157eb4fb_result_delayed_result_delayed_u0<=1'h0;
else reg_157eb4fb_result_delayed_result_delayed_u0<=reg_157eb4fb_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4a382354_result_delayed_u0<=1'h0;
else reg_4a382354_result_delayed_u0<=reg_4a382354_u0;
end
assign and_u1765_u0=and_u1759_u0&and_u1767_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0e249eb7_result_delayed_u0<=1'h0;
else reg_0e249eb7_result_delayed_u0<=reg_0e249eb7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1bd6ae3f_result_delayed_result_delayed_u0<=1'h0;
else reg_1bd6ae3f_result_delayed_result_delayed_u0<=reg_1bd6ae3f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2c6d2fd0_u0<=1'h0;
else reg_2c6d2fd0_u0<=reg_216d1570_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0dc8a158_result_delayed_u0<=1'h0;
else reg_0dc8a158_result_delayed_u0<=reg_0dc8a158_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_216d1570_result_delayed_result_delayed_u0<=1'h0;
else reg_216d1570_result_delayed_result_delayed_u0<=reg_216d1570_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_72f7e7fe_result_delayed_u0<=1'h0;
else reg_72f7e7fe_result_delayed_u0<=reg_72f7e7fe_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2ab2a055_result_delayed_u0<=1'h0;
else reg_2ab2a055_result_delayed_u0<=reg_2ab2a055_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2b4cee92_result_delayed_u0<=1'h0;
else reg_2b4cee92_result_delayed_u0<=reg_2b4cee92_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_16db469f_result_delayed_u0<=1'h0;
else reg_16db469f_result_delayed_u0<=reg_16db469f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4bc0004f_result_delayed_u0<=1'h0;
else reg_4bc0004f_result_delayed_u0<=reg_4bc0004f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2e9b949b_result_delayed_u0<=1'h0;
else reg_2e9b949b_result_delayed_u0<=reg_2e9b949b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_07979748_result_delayed_result_delayed_u0<=1'h0;
else reg_07979748_result_delayed_result_delayed_u0<=reg_07979748_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4bfc6bcc_result_delayed_result_delayed_u0<=1'h0;
else reg_4bfc6bcc_result_delayed_result_delayed_u0<=reg_4bfc6bcc_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_297e0532_result_delayed_u0<=1'h0;
else reg_297e0532_result_delayed_u0<=reg_297e0532_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1bd6ae3f_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_1bd6ae3f_result_delayed_result_delayed_result_delayed_u0<=reg_1bd6ae3f_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_776a1f94_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_776a1f94_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_776a1f94_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_74845d78_result_delayed_u0<=1'h0;
else reg_74845d78_result_delayed_u0<=reg_74845d78_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_247a1111_result_delayed_u0<=1'h0;
else reg_247a1111_result_delayed_u0<=reg_247a1111_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_30bea5e3_result_delayed_result_delayed_u0<=1'h0;
else reg_30bea5e3_result_delayed_result_delayed_u0<=reg_30bea5e3_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_170037b2_result_delayed_result_delayed_u0<=1'h0;
else reg_170037b2_result_delayed_result_delayed_u0<=reg_170037b2_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_319759b9_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_319759b9_result_delayed_result_delayed_result_delayed_u0<=reg_319759b9_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_63d04af9_result_delayed_result_delayed_u0<=1'h0;
else reg_63d04af9_result_delayed_result_delayed_u0<=reg_63d04af9_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6ee280fb_result_delayed_u0<=1'h0;
else reg_6ee280fb_result_delayed_u0<=reg_6ee280fb_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3771f97a_result_delayed_u0<=1'h0;
else reg_3771f97a_result_delayed_u0<=reg_3771f97a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_44a091fd_result_delayed_u0<=1'h0;
else reg_44a091fd_result_delayed_u0<=reg_44a091fd_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5c0a547e_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_5c0a547e_result_delayed_result_delayed_result_delayed_u0<=reg_5c0a547e_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a591648_result_delayed_result_delayed_u0<=1'h0;
else reg_7a591648_result_delayed_result_delayed_u0<=reg_7a591648_result_delayed_u0;
end
assign or_u483_u0=and_u1766_u0|and_u1765_u0;
assign or_u484_u0=and_delayed_result_delayed_result_delayed_u2|or_u481_u0;
assign mux_u181_u0=(and_u1766_u0)?1'h1:mux_u180;
assign or_u485_u0=and_u1766_u0|or_u482_u0;
assign and_u1766_u0=and_u1758_u0&and_u1769_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u118<=1'h0;
else and_delayed_u118<=and_u1766_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_result_delayed_u9<=1'h0;
else and_delayed_result_delayed_u9<=and_delayed_u118;
end
assign and_u1767_u0=and_u1757_u0&and_u1769_u0;
assign or_u486_u0=and_u1766_u0|and_u1765_u0;
assign mux_u182_u0=(and_u1766_u0)?32'h2:32'h200;
assign or_u487_u0=and_u1766_u0|and_u1765_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_result_delayed_result_delayed_u2<=1'h0;
else and_delayed_result_delayed_result_delayed_u2<=and_delayed_result_delayed_u9;
end
assign or_u488_u0=and_u1766_u0|and_u1765_u0;
assign and_u1768_u0=and_u1756_u0&and_u1754_u0;
assign or_u489_u0=and_delayed_u119_u0|or_u484_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u119_u0<=1'h0;
else and_delayed_u119_u0<=and_u1768_u0;
end
assign and_u1769_u0=and_u1755_u0&and_u1754_u0;
assign equals_u94_a_signed={31'b0, port_0712fa18_};
assign equals_u94_b_signed=32'h1;
assign equals_u94=equals_u94_a_signed==equals_u94_b_signed;
assign and_u1770_u0=and_u1754_u0&equals_u94;
assign and_u1771_u0=and_u1754_u0&not_u350_u0;
assign not_u350_u0=~equals_u94;
assign and_u1772_u0=and_u1786_u0&not_u351_u0;
assign and_u1773_u0=and_u1786_u0&port_35218c17_;
assign not_u351_u0=~port_35218c17_;
assign lessThan_u39_a_signed=port_5ff18c4c_;
assign lessThan_u39_b_signed=port_4c4a747e_;
assign lessThan_u39=lessThan_u39_a_signed<lessThan_u39_b_signed;
assign not_u352_u0=~lessThan_u39;
assign and_u1774_u0=and_u1784_u0&not_u352_u0;
assign and_u1775_u0=and_u1784_u0&lessThan_u39;
assign not_u353_u0=~port_6b386c73_;
assign and_u1776_u0=and_u1781_u0&port_6b386c73_;
assign and_u1777_u0=and_u1781_u0&not_u353_u0;
assign add=port_5ff18c4c_+32'h0;
assign and_u1778_u0=and_u1780_u0&port_27356da8_;
assign simplePinWrite_u318=16'h1&{16{1'h1}};
assign simplePinWrite_u319=port_72850e0c_;
assign simplePinWrite_u320=and_u1780_u0&{1{and_u1780_u0}};
assign add_u68=port_5ff18c4c_+32'h1;
always @(posedge CLK)
begin
if (and_u1780_u0)
syncEnable_u180<=port_72850e0c_;
end
assign mux_u183_u0=(and_delayed_u120_u0)?syncEnable_u181_u0:syncEnable_u180;
assign and_u1779_u0=and_u1777_u0&and_u1781_u0;
assign and_u1780_u0=and_u1776_u0&and_u1781_u0;
always @(posedge CLK)
begin
if (and_u1781_u0)
syncEnable_u181_u0<=mux_u195_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u120_u0<=1'h0;
else and_delayed_u120_u0<=and_u1779_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u121_u0<=1'h0;
else and_delayed_u121_u0<=and_u1780_u0;
end
always @(posedge CLK)
begin
if (and_u1784_u0)
syncEnable_u182_u0<=mux_u194_u0;
end
assign mux_u184_u0=(reg_645b9fd5_u0)?syncEnable_u183_u0:mux_u183_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4dcef723_u0<=1'h0;
else reg_4dcef723_u0<=and_u1781_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_645b9fd5_u0<=1'h0;
else reg_645b9fd5_u0<=and_u1782_u0;
end
assign and_u1781_u0=and_u1775_u0&and_u1784_u0;
always @(posedge CLK)
begin
if (and_u1784_u0)
syncEnable_u183_u0<=mux_u195_u0;
end
assign and_u1782_u0=and_u1774_u0&and_u1784_u0;
assign mux_u185_u0=(reg_645b9fd5_u0)?32'h0:syncEnable_u182_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1a01de45_u0<=1'h0;
else reg_1a01de45_u0<=and_u1783_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_535070be_u0<=1'h0;
else reg_535070be_u0<=and_u1784_u0;
end
always @(posedge CLK)
begin
if (and_u1786_u0)
syncEnable_u184_u0<=mux_u194_u0;
end
assign and_u1783_u0=and_u1772_u0&and_u1786_u0;
assign and_u1784_u0=and_u1773_u0&and_u1786_u0;
assign mux_u186_u0=(reg_535070be_u0)?mux_u185_u0:syncEnable_u184_u0;
assign mux_u187_u0=(reg_535070be_u0)?mux_u184_u0:syncEnable_u185_u0;
always @(posedge CLK)
begin
if (and_u1786_u0)
syncEnable_u185_u0<=mux_u195_u0;
end
assign mux_u188_u0=(and_delayed_u122_u0)?mux_u187_u0:syncEnable_u187_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5039c73f_u0<=1'h0;
else reg_5039c73f_u0<=and_u1785_u0;
end
assign and_u1785_u0=and_u1771_u0&and_u1754_u0;
always @(posedge CLK)
begin
if (and_u1754_u0)
syncEnable_u186_u0<=mux_u194_u0;
end
assign and_u1786_u0=and_u1770_u0&and_u1754_u0;
assign mux_u189_u0=(and_delayed_u122_u0)?mux_u186_u0:syncEnable_u186_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u122_u0<=1'h0;
else and_delayed_u122_u0<=and_u1786_u0;
end
always @(posedge CLK)
begin
if (and_u1754_u0)
syncEnable_u187_u0<=mux_u195_u0;
end
assign mux_u190_u0=(or_u485_u0)?mux_u181_u0:1'h0;
assign or_u490_u0=or_u485_u0|and_u1782_u0;
assign latch_4d9bcb18_out=(block_GO_delayed_u6)?mux_u188_u0:latch_4d9bcb18_reg;
always @(posedge CLK)
begin
if (block_GO_delayed_u6)
latch_4d9bcb18_reg<=mux_u188_u0;
end
assign or_u491_u0=or_u483_u0|and_u1780_u0;
assign mux_u191_u0=(or_u483_u0)?32'h0:add_u68;
assign latch_1e7607d8_out=(block_GO_delayed_u6)?mux_u189_u0:latch_1e7607d8_reg;
always @(posedge CLK)
begin
if (block_GO_delayed_u6)
latch_1e7607d8_reg<=mux_u189_u0;
end
assign or_u492_u0=or_u487_u0|and_u1782_u0;
assign mux_u192_u0=(or_u487_u0)?1'h1:1'h0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
block_GO_delayed_u6<=1'h0;
else block_GO_delayed_u6<=and_u1754_u0;
end
assign or_u493_u0=or_u486_u0|and_u1782_u0;
assign mux_u193_u0=(or_u486_u0)?{22'b0, mux_u182_u0[9], 7'b0, mux_u182_u0[1], 1'b0}:32'hffffffff;
assign mux_u194_u0=(reg_36b6d836_result_delayed_u0)?32'h0:fbReg_temp_fsmOldState_resized_HH1_xy_3_u0;
assign or_u494_u0=reg_36b6d836_result_delayed_u0|loopControl_u3;
always @(posedge CLK)
begin
if (or_u489_u0)
fbReg_temp_fsmOldState_resized_HH1_xy_3_u0<=latch_1e7607d8_out;
end
always @(posedge CLK or posedge syncEnable_u188_u0)
begin
if (syncEnable_u188_u0)
loopControl_u3<=1'h0;
else loopControl_u3<=or_u489_u0;
end
assign mux_u195_u0=(reg_36b6d836_result_delayed_u0)?16'h0:fbReg_Out1Portvalue_u0;
always @(posedge CLK)
begin
if (reg_36b6d836_result_delayed_u0)
syncEnable_u188_u0<=RESET;
end
always @(posedge CLK)
begin
if (or_u489_u0)
fbReg_Out1Portvalue_u0<=latch_4d9bcb18_out;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_36b6d836_u0<=1'h0;
else reg_36b6d836_u0<=GO;
end
assign or_u495_u0=GO|or_u491_u0;
assign mux_u196_u0=(GO)?32'h0:mux_u191_u0;
assign or_u496_u0=GO|or_u488_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_36b6d836_result_delayed_u0<=1'h0;
else reg_36b6d836_result_delayed_u0<=reg_36b6d836_u0;
end
assign or_u497_u0=GO|or_u493_u0;
assign mux_u197_u0=(GO)?32'hffffffff:mux_u193_u0;
assign or_u498_u0=GO|or_u490_u0;
assign mux_u198_u0=(GO)?1'h0:mux_u190_u0;
assign or_u499_u0=GO|or_u492_u0;
assign mux_u199_u0=(GO)?1'h0:mux_u192_u0;
assign RESULT=or_u496_u0;
assign RESULT_u1083=32'h0;
assign RESULT_u1084=or_u498_u0;
assign RESULT_u1085=mux_u198_u0;
assign RESULT_u1086=or_u495_u0;
assign RESULT_u1087=mux_u196_u0;
assign RESULT_u1088=or_u497_u0;
assign RESULT_u1089=mux_u197_u0;
assign RESULT_u1090=or_u499_u0;
assign RESULT_u1091=mux_u199_u0;
assign RESULT_u1092=and_u1780_u0;
assign RESULT_u1093=add;
assign RESULT_u1094=3'h1;
assign RESULT_u1095=simplePinWrite;
assign RESULT_u1096=simplePinWrite_u318;
assign RESULT_u1097=simplePinWrite_u316;
assign RESULT_u1098=simplePinWrite_u320;
assign RESULT_u1099=simplePinWrite_u317;
assign RESULT_u1100=simplePinWrite_u319;
assign DONE=1'h0;
endmodule



module resized_HH1_xy_structuralmemory_4abb499d_(CLK_u9, bus_20b8f358_, bus_233a1a3f_, bus_2226f9ce_, bus_7cf55b9c_, bus_5deb4f38_, bus_2319feae_, bus_7b7cec0a_, bus_0ec3b904_);
input		CLK_u9;
input		bus_20b8f358_;
input	[31:0]	bus_233a1a3f_;
input	[2:0]	bus_2226f9ce_;
input		bus_7cf55b9c_;
input		bus_5deb4f38_;
input	[15:0]	bus_2319feae_;
output	[15:0]	bus_7b7cec0a_;
output		bus_0ec3b904_;
reg		logicalMem_5a9b60d1_we_delay0_u0=1'h0;
wire	[15:0]	bus_4ea56e93_;
wire		not_5bbc05c8_u0;
wire		and_3ce245b7_u0;
wire		or_733d2261_u0;
wire		or_0bfcd463_u0;
always @(posedge CLK_u9 or posedge bus_20b8f358_)
begin
if (bus_20b8f358_)
logicalMem_5a9b60d1_we_delay0_u0<=1'h0;
else logicalMem_5a9b60d1_we_delay0_u0<=bus_5deb4f38_;
end
assign bus_7b7cec0a_=bus_4ea56e93_;
assign bus_0ec3b904_=or_733d2261_u0;
resized_HH1_xy_forge_memory_512x16_18 resized_HH1_xy_forge_memory_512x16_18_instance1(.CLK(CLK_u9), 
  .EN(or_0bfcd463_u0), .WE(bus_5deb4f38_), .ADDR(bus_233a1a3f_), .DIN(bus_2319feae_), 
  .DOUT(bus_4ea56e93_), .DONE());
assign not_5bbc05c8_u0=~bus_5deb4f38_;
assign and_3ce245b7_u0=bus_7cf55b9c_&not_5bbc05c8_u0;
assign or_733d2261_u0=and_3ce245b7_u0|logicalMem_5a9b60d1_we_delay0_u0;
assign or_0bfcd463_u0=bus_7cf55b9c_|bus_5deb4f38_;
endmodule



module resized_HH1_xy_reset(CLK, RESET, GO, RESULT, RESULT_u1101, RESULT_u1102, RESULT_u1103, DONE);
input		CLK;
input		RESET;
input		GO;
output		RESULT;
output	[15:0]	RESULT_u1101;
output		RESULT_u1102;
output	[15:0]	RESULT_u1103;
output		DONE;
reg		reg_571be4a7_u0=1'h0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_571be4a7_u0<=1'h0;
else reg_571be4a7_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u1101=16'h1;
assign RESULT_u1102=GO;
assign RESULT_u1103=16'h0;
assign DONE=reg_571be4a7_u0;
endmodule



module resized_HH1_xy_globalreset_physical_35a1308a_(bus_61966029_, bus_12c51121_, bus_1d017b90_);
input		bus_61966029_;
input		bus_12c51121_;
output		bus_1d017b90_;
wire		or_647926ab_u0;
reg		glitch_u33=1'h0;
reg		sample_u33=1'h0;
reg		cross_u33=1'h0;
reg		final_u33=1'h1;
wire		not_6439c7b2_u0;
wire		and_7e695774_u0;
assign bus_1d017b90_=or_647926ab_u0;
assign or_647926ab_u0=bus_12c51121_|final_u33;
always @(posedge bus_61966029_)
begin
glitch_u33<=cross_u33;
end
always @(posedge bus_61966029_)
begin
sample_u33<=1'h1;
end
always @(posedge bus_61966029_)
begin
cross_u33<=sample_u33;
end
always @(posedge bus_61966029_)
begin
final_u33<=not_6439c7b2_u0;
end
assign not_6439c7b2_u0=~and_7e695774_u0;
assign and_7e695774_u0=cross_u33&glitch_u33;
endmodule



module resized_HH1_xy_endianswapper_25188211_(endianswapper_25188211_in, endianswapper_25188211_out);
input	[31:0]	endianswapper_25188211_in;
output	[31:0]	endianswapper_25188211_out;
assign endianswapper_25188211_out=endianswapper_25188211_in;
endmodule



module resized_HH1_xy_endianswapper_7e80f5bd_(endianswapper_7e80f5bd_in, endianswapper_7e80f5bd_out);
input	[31:0]	endianswapper_7e80f5bd_in;
output	[31:0]	endianswapper_7e80f5bd_out;
assign endianswapper_7e80f5bd_out=endianswapper_7e80f5bd_in;
endmodule



module resized_HH1_xy_stateVar_Out1TokenIndex(bus_4d2a4e2c_, bus_65b626e0_, bus_4a4819b0_, bus_01d9d88c_, bus_7fd1c7f0_);
input		bus_4d2a4e2c_;
input		bus_65b626e0_;
input		bus_4a4819b0_;
input	[31:0]	bus_01d9d88c_;
output	[31:0]	bus_7fd1c7f0_;
reg	[31:0]	stateVar_Out1TokenIndex_u0=32'h0;
wire	[31:0]	endianswapper_25188211_out;
wire	[31:0]	endianswapper_7e80f5bd_out;
always @(posedge bus_4d2a4e2c_ or posedge bus_65b626e0_)
begin
if (bus_65b626e0_)
stateVar_Out1TokenIndex_u0<=32'h0;
else if (bus_4a4819b0_)
stateVar_Out1TokenIndex_u0<=endianswapper_25188211_out;
end
assign bus_7fd1c7f0_=endianswapper_7e80f5bd_out;
resized_HH1_xy_endianswapper_25188211_ resized_HH1_xy_endianswapper_25188211__1(.endianswapper_25188211_in(bus_01d9d88c_), 
  .endianswapper_25188211_out(endianswapper_25188211_out));
resized_HH1_xy_endianswapper_7e80f5bd_ resized_HH1_xy_endianswapper_7e80f5bd__1(.endianswapper_7e80f5bd_in(stateVar_Out1TokenIndex_u0), 
  .endianswapper_7e80f5bd_out(endianswapper_7e80f5bd_out));
endmodule



module resized_HH1_xy_endianswapper_601849ef_(endianswapper_601849ef_in, endianswapper_601849ef_out);
input	[15:0]	endianswapper_601849ef_in;
output	[15:0]	endianswapper_601849ef_out;
assign endianswapper_601849ef_out=endianswapper_601849ef_in;
endmodule



module resized_HH1_xy_endianswapper_4fde4273_(endianswapper_4fde4273_in, endianswapper_4fde4273_out);
input	[15:0]	endianswapper_4fde4273_in;
output	[15:0]	endianswapper_4fde4273_out;
assign endianswapper_4fde4273_out=endianswapper_4fde4273_in;
endmodule



module resized_HH1_xy_stateVar_rowRepeated(bus_19552c76_, bus_590dd011_, bus_52fff2e1_, bus_55439b52_, bus_6a21e216_, bus_0bb2ece1_, bus_46857e3b_);
input		bus_19552c76_;
input		bus_590dd011_;
input		bus_52fff2e1_;
input	[15:0]	bus_55439b52_;
input		bus_6a21e216_;
input	[15:0]	bus_0bb2ece1_;
output	[15:0]	bus_46857e3b_;
wire	[15:0]	endianswapper_601849ef_out;
wire	[15:0]	mux_3b26358e_u0;
reg	[15:0]	stateVar_rowRepeated_u0=16'h1;
wire		or_307cbd16_u0;
wire	[15:0]	endianswapper_4fde4273_out;
resized_HH1_xy_endianswapper_601849ef_ resized_HH1_xy_endianswapper_601849ef__1(.endianswapper_601849ef_in(stateVar_rowRepeated_u0), 
  .endianswapper_601849ef_out(endianswapper_601849ef_out));
assign mux_3b26358e_u0=(bus_52fff2e1_)?bus_55439b52_:16'h1;
always @(posedge bus_19552c76_ or posedge bus_590dd011_)
begin
if (bus_590dd011_)
stateVar_rowRepeated_u0<=16'h1;
else if (or_307cbd16_u0)
stateVar_rowRepeated_u0<=endianswapper_4fde4273_out;
end
assign bus_46857e3b_=endianswapper_601849ef_out;
assign or_307cbd16_u0=bus_52fff2e1_|bus_6a21e216_;
resized_HH1_xy_endianswapper_4fde4273_ resized_HH1_xy_endianswapper_4fde4273__1(.endianswapper_4fde4273_in(mux_3b26358e_u0), 
  .endianswapper_4fde4273_out(endianswapper_4fde4273_out));
endmodule



module resized_HH1_xy_consumeRow(CLK, RESET, GO, port_531ffb68_, port_402540c6_, port_0d7ca19e_, port_2e5e0079_, RESULT, RESULT_u1104, RESULT_u1105, RESULT_u1106, RESULT_u1107, RESULT_u1108, RESULT_u1109, RESULT_u1110, RESULT_u1111, RESULT_u1112, RESULT_u1113, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_531ffb68_;
input		port_402540c6_;
input		port_0d7ca19e_;
input	[15:0]	port_2e5e0079_;
output		RESULT;
output	[15:0]	RESULT_u1104;
output		RESULT_u1105;
output	[31:0]	RESULT_u1106;
output	[15:0]	RESULT_u1107;
output	[2:0]	RESULT_u1108;
output		RESULT_u1109;
output	[31:0]	RESULT_u1110;
output	[15:0]	RESULT_u1111;
output	[2:0]	RESULT_u1112;
output		RESULT_u1113;
output		DONE;
wire		simplePinWrite;
wire	[31:0]	add;
wire	[31:0]	add_u69;
reg		reg_6112dc10_u0=1'h0;
wire		and_u1787_u0;
wire		or_u500_u0;
wire	[15:0]	add_u70;
reg	[15:0]	syncEnable_u189=16'h0;
reg		reg_33a16981_u0=1'h0;
wire		and_u1788_u0;
wire		and_u1789_u0;
wire signed	[16:0]	lessThanEqualTo_a_signed;
wire signed	[16:0]	lessThanEqualTo_b_signed;
wire		lessThanEqualTo;
wire		and_u1790_u0;
wire		and_u1791_u0;
wire		not_u354_u0;
wire		or_u501_u0;
reg	[15:0]	latch_79398a8d_reg=16'h0;
wire	[15:0]	latch_79398a8d_out;
wire	[15:0]	mux_u200;
wire	[15:0]	add_u71;
wire		lessThanEqualTo_u0;
wire signed	[16:0]	lessThanEqualTo_u0_a_signed;
wire signed	[16:0]	lessThanEqualTo_u0_b_signed;
wire		and_u1792_u0;
wire		not_u355_u0;
wire		and_u1793_u0;
reg		reg_5be3984a_u0=1'h0;
wire		and_u1794_u0;
wire	[15:0]	subtract;
wire	[31:0]	add_u72;
wire		or_u502_u0;
wire		and_u1795_u0;
reg		reg_70cfdd52_u0=1'h0;
wire	[15:0]	add_u73;
reg	[15:0]	syncEnable_u190_u0=16'h0;
wire		and_u1796_u0;
wire		or_u503_u0;
wire	[15:0]	mux_u201_u0;
wire	[15:0]	latch_5ee2d6fa_out;
reg	[15:0]	latch_5ee2d6fa_reg=16'h0;
reg	[15:0]	syncEnable_u191_u0=16'h0;
reg		reg_79389cc5_u0=1'h0;
assign simplePinWrite=GO&{1{GO}};
assign add={15'b0, port_531ffb68_, 1'b0}+{mux_u200[15], mux_u200[15], mux_u200[15], mux_u200[15], mux_u200[15], mux_u200[15], mux_u200[15], mux_u200[15], mux_u200[15], mux_u200[15], mux_u200[15], mux_u200[15], mux_u200[15], mux_u200[15], mux_u200[15], mux_u200[15], mux_u200};
assign add_u69={add[18], add[18], add[18], add[18], add[18], add[18], add[18], add[18], add[18], add[18], add[18], add[18], add[18], add[18:0]}+32'h0;
always @(posedge CLK or posedge and_u1789_u0 or posedge or_u500_u0)
begin
if (or_u500_u0)
reg_6112dc10_u0<=1'h0;
else if (and_u1789_u0)
reg_6112dc10_u0<=1'h1;
else reg_6112dc10_u0<=reg_6112dc10_u0;
end
assign and_u1787_u0=reg_6112dc10_u0&port_0d7ca19e_;
assign or_u500_u0=and_u1787_u0|RESET;
assign add_u70=mux_u200+16'h1;
always @(posedge CLK)
begin
if (and_u1789_u0)
syncEnable_u189<=add_u70;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_33a16981_u0<=1'h0;
else reg_33a16981_u0<=and_u1789_u0;
end
assign and_u1788_u0=and_u1791_u0&or_u501_u0;
assign and_u1789_u0=and_u1790_u0&or_u501_u0;
assign lessThanEqualTo_a_signed={mux_u200[15], mux_u200};
assign lessThanEqualTo_b_signed=17'h1;
assign lessThanEqualTo=lessThanEqualTo_a_signed<=lessThanEqualTo_b_signed;
assign and_u1790_u0=or_u501_u0&lessThanEqualTo;
assign and_u1791_u0=or_u501_u0&not_u354_u0;
assign not_u354_u0=~lessThanEqualTo;
assign or_u501_u0=reg_33a16981_u0|GO;
always @(posedge CLK)
begin
if (GO)
latch_79398a8d_reg<=port_2e5e0079_;
end
assign latch_79398a8d_out=(GO)?port_2e5e0079_:latch_79398a8d_reg;
assign mux_u200=(reg_33a16981_u0)?syncEnable_u189:16'h0;
assign add_u71=port_531ffb68_+16'h1;
assign lessThanEqualTo_u0_a_signed={mux_u201_u0[15], mux_u201_u0};
assign lessThanEqualTo_u0_b_signed=17'h2;
assign lessThanEqualTo_u0=lessThanEqualTo_u0_a_signed<=lessThanEqualTo_u0_b_signed;
assign and_u1792_u0=or_u503_u0&lessThanEqualTo_u0;
assign not_u355_u0=~lessThanEqualTo_u0;
assign and_u1793_u0=or_u503_u0&not_u355_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5be3984a_u0<=1'h0;
else reg_5be3984a_u0<=and_u1796_u0;
end
assign and_u1794_u0=and_u1793_u0&or_u503_u0;
assign subtract=mux_u201_u0-16'h1;
assign add_u72={subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract}+32'h0;
assign or_u502_u0=and_u1795_u0|RESET;
assign and_u1795_u0=reg_70cfdd52_u0&port_402540c6_;
always @(posedge CLK or posedge and_u1796_u0 or posedge or_u502_u0)
begin
if (or_u502_u0)
reg_70cfdd52_u0<=1'h0;
else if (and_u1796_u0)
reg_70cfdd52_u0<=1'h1;
else reg_70cfdd52_u0<=reg_70cfdd52_u0;
end
assign add_u73=mux_u201_u0+16'h1;
always @(posedge CLK)
begin
if (and_u1796_u0)
syncEnable_u190_u0<=add_u73;
end
assign and_u1796_u0=and_u1792_u0&or_u503_u0;
assign or_u503_u0=GO|reg_5be3984a_u0;
assign mux_u201_u0=(GO)?16'h1:syncEnable_u190_u0;
assign latch_5ee2d6fa_out=(GO)?port_2e5e0079_:latch_5ee2d6fa_reg;
always @(posedge CLK)
begin
if (GO)
latch_5ee2d6fa_reg<=port_2e5e0079_;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u191_u0<=add_u71;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_79389cc5_u0<=1'h0;
else reg_79389cc5_u0<=and_u1788_u0;
end
assign RESULT=and_u1788_u0;
assign RESULT_u1104=syncEnable_u191_u0;
assign RESULT_u1105=and_u1796_u0;
assign RESULT_u1106=add_u72;
assign RESULT_u1107=latch_5ee2d6fa_out;
assign RESULT_u1108=3'h1;
assign RESULT_u1109=and_u1789_u0;
assign RESULT_u1110=add_u69;
assign RESULT_u1111=latch_79398a8d_out;
assign RESULT_u1112=3'h1;
assign RESULT_u1113=simplePinWrite;
assign DONE=reg_79389cc5_u0;
endmodule


