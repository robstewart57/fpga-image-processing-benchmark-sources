// __  ___ __ ___  _ __   ___  ___ 
// \ \/ / '__/ _ \| '_ \ / _ \/ __|
//  >  <| | | (_) | | | | (_) \__ \
// /_/\_\_|  \___/|_| |_|\___/|___/
// 
// Xronos synthesizer version
// Run date: Thu 2 Nov 2017 13:59:32 +0000
// 

module resized_LH2_xy(In1_ACK, In1_COUNT, Out1_DATA, Out1_SEND, Out1_COUNT, Out1_ACK, CLK, In1_DATA, RESET, In1_SEND, Out1_RDY);
output		In1_ACK;
input	[15:0]	In1_COUNT;
output	[15:0]	Out1_DATA;
wire		reset_done;
output		Out1_SEND;
output	[15:0]	Out1_COUNT;
input		Out1_ACK;
input		CLK;
wire		consumeRow_go;
input	[15:0]	In1_DATA;
wire		reset_go;
input		RESET;
input		In1_SEND;
input		Out1_RDY;
wire		repeatRowExpanded_go;
wire		repeatRowExpanded_done;
wire		consumeRow_done;
wire		bus_4a33a20e_;
wire	[15:0]	bus_703c1161_;
wire		bus_7fd3fe0c_;
wire		bus_5895103d_;
wire	[31:0]	bus_5bffa9c0_;
wire	[31:0]	bus_7281aa61_;
wire	[31:0]	bus_3b01d7ce_;
wire	[2:0]	repeatRowExpanded_u39;
wire		repeatRowExpanded_u33;
wire		repeatRowExpanded_u37;
wire		repeatRowExpanded;
wire	[2:0]	repeatRowExpanded_u36;
wire	[31:0]	repeatRowExpanded_u38;
wire	[15:0]	repeatRowExpanded_u35;
wire		resized_LH2_xy_repeatRowExpanded_instance_DONE;
wire	[15:0]	repeatRowExpanded_u32;
wire	[31:0]	repeatRowExpanded_u34;
wire		bus_0e8f38dd_;
wire	[31:0]	bus_706839bc_;
wire	[2:0]	bus_551a77e4_;
wire	[15:0]	bus_01a9e6ce_;
wire		bus_1bceed37_;
wire		bus_768c4387_;
wire		bus_1307238a_;
wire	[15:0]	bus_4bbace21_;
wire	[31:0]	scheduler_u309;
wire		scheduler_u313;
wire		scheduler_u308;
wire		scheduler_u300;
wire		scheduler_u302;
wire		scheduler_u311;
wire		scheduler_u307;
wire		resized_LH2_xy_scheduler_instance_DONE;
wire	[31:0]	scheduler_u303;
wire		scheduler_u306;
wire	[2:0]	scheduler_u310;
wire		scheduler_u314;
wire		scheduler_u304;
wire		scheduler;
wire	[15:0]	scheduler_u312;
wire		scheduler_u315;
wire	[31:0]	scheduler_u305;
wire	[31:0]	scheduler_u299;
wire		scheduler_u301;
wire	[15:0]	scheduler_u316;
wire	[15:0]	bus_45cec17e_;
wire	[15:0]	bus_2b80c1a2_;
wire		bus_2bfcb357_;
wire		resized_LH2_xy_reset_instance_DONE;
wire	[15:0]	reset_u12;
wire		reset_u13;
wire	[15:0]	reset_u14;
wire		reset;
wire		bus_7aafd725_;
wire		bus_112f0657_;
wire		consumeRow;
wire	[15:0]	consumeRow_u40;
wire	[15:0]	consumeRow_u47;
wire		consumeRow_u49;
wire	[2:0]	consumeRow_u44;
wire		consumeRow_u45;
wire	[2:0]	consumeRow_u48;
wire		resized_LH2_xy_consumeRow_instance_DONE;
wire	[15:0]	consumeRow_u43;
wire	[31:0]	consumeRow_u42;
wire	[31:0]	consumeRow_u46;
wire		consumeRow_u41;
wire		bus_2a450b51_;
wire	[15:0]	bus_0f871660_;
wire		bus_55b75661_;
wire		bus_52d26b67_;
wire	[15:0]	bus_4686658d_;
wire		bus_736af7eb_;
wire		bus_04f85a99_;
wire		bus_4687e307_;
wire		bus_307decb9_;
wire		bus_13df4b68_;
wire	[2:0]	bus_50563d51_;
wire	[31:0]	bus_05401935_;
wire	[15:0]	bus_180d93a2_;
assign In1_ACK=consumeRow_u49;
assign Out1_DATA=scheduler_u316;
assign reset_done=bus_7fd3fe0c_;
assign Out1_SEND=scheduler_u311;
assign Out1_COUNT=scheduler_u312;
assign consumeRow_go=scheduler_u314;
assign reset_go=scheduler_u315;
assign repeatRowExpanded_go=scheduler_u313;
assign repeatRowExpanded_done=bus_7aafd725_;
assign consumeRow_done=bus_5895103d_;
resized_LH2_xy_Kicker_45 resized_LH2_xy_Kicker_45_1(.CLK(CLK), .RESET(bus_112f0657_), 
  .bus_4a33a20e_(bus_4a33a20e_));
resized_LH2_xy_stateVar_x resized_LH2_xy_stateVar_x_1(.bus_49987487_(CLK), .bus_5d8644af_(bus_112f0657_), 
  .bus_551d1965_(consumeRow), .bus_30e7f77b_(consumeRow_u40), .bus_75dc4e7a_(reset_u13), 
  .bus_7e3885be_(16'h0), .bus_703c1161_(bus_703c1161_));
assign bus_7fd3fe0c_=resized_LH2_xy_reset_instance_DONE&{1{resized_LH2_xy_reset_instance_DONE}};
assign bus_5895103d_=resized_LH2_xy_consumeRow_instance_DONE&{1{resized_LH2_xy_consumeRow_instance_DONE}};
resized_LH2_xy_stateVar_fsmOldState_resized_LH2_xy resized_LH2_xy_stateVar_fsmOldState_resized_LH2_xy_1(.bus_38a242af_(CLK), 
  .bus_3a6e3652_(bus_112f0657_), .bus_54189c3e_(scheduler), .bus_35927e1c_(32'h0), 
  .bus_5bffa9c0_(bus_5bffa9c0_));
resized_LH2_xy_stateVar_Out1MaxTokenIndex resized_LH2_xy_stateVar_Out1MaxTokenIndex_1(.bus_7d661b62_(CLK), 
  .bus_26c83530_(bus_112f0657_), .bus_691cf5a3_(scheduler_u304), .bus_43ea8ee1_(scheduler_u305), 
  .bus_7281aa61_(bus_7281aa61_));
resized_LH2_xy_stateVar_Out1TokenIndex resized_LH2_xy_stateVar_Out1TokenIndex_1(.bus_71cf89b8_(CLK), 
  .bus_1502dffb_(bus_112f0657_), .bus_2791719c_(scheduler_u302), .bus_29e05130_(scheduler_u303), 
  .bus_3b01d7ce_(bus_3b01d7ce_));
resized_LH2_xy_repeatRowExpanded resized_LH2_xy_repeatRowExpanded_instance(.CLK(CLK), 
  .RESET(bus_112f0657_), .GO(repeatRowExpanded_go), .port_5bf0021c_(bus_45cec17e_), 
  .port_2dd6a8c5_(bus_307decb9_), .port_3f45710a_(bus_768c4387_), .port_047547ec_(bus_4bbace21_), 
  .DONE(resized_LH2_xy_repeatRowExpanded_instance_DONE), .RESULT(repeatRowExpanded), 
  .RESULT_u2111(repeatRowExpanded_u32), .RESULT_u2112(repeatRowExpanded_u33), 
  .RESULT_u2113(repeatRowExpanded_u34), .RESULT_u2114(repeatRowExpanded_u35), 
  .RESULT_u2115(repeatRowExpanded_u36), .RESULT_u2116(repeatRowExpanded_u37), 
  .RESULT_u2117(repeatRowExpanded_u38), .RESULT_u2118(repeatRowExpanded_u39));
resized_LH2_xy_simplememoryreferee_53c3fe95_ resized_LH2_xy_simplememoryreferee_53c3fe95__1(.bus_329d11ec_(CLK), 
  .bus_6055eb84_(bus_112f0657_), .bus_23b69ded_(bus_2bfcb357_), .bus_0d07a037_(bus_2b80c1a2_), 
  .bus_42291ec9_(consumeRow_u41), .bus_4d695e2f_(consumeRow_u43), .bus_6f653eab_(consumeRow_u42), 
  .bus_7bc2b5e6_(3'h1), .bus_277138ad_(repeatRowExpanded_u37), .bus_278380fd_(repeatRowExpanded_u38), 
  .bus_34fe08d6_(3'h1), .bus_01a9e6ce_(bus_01a9e6ce_), .bus_706839bc_(bus_706839bc_), 
  .bus_0e8f38dd_(bus_0e8f38dd_), .bus_1307238a_(bus_1307238a_), .bus_551a77e4_(bus_551a77e4_), 
  .bus_1bceed37_(bus_1bceed37_), .bus_4bbace21_(bus_4bbace21_), .bus_768c4387_(bus_768c4387_));
resized_LH2_xy_scheduler resized_LH2_xy_scheduler_instance(.CLK(CLK), .RESET(bus_112f0657_), 
  .GO(bus_4a33a20e_), .port_3b0b1e1a_(32'h0), .port_5b3d11e3_(bus_2a450b51_), .port_5aad7090_(bus_3b01d7ce_), 
  .port_598dd3c9_(bus_7281aa61_), .port_02986e5e_(bus_52d26b67_), .port_177051de_(bus_703c1161_), 
  .port_386b1b7a_(bus_45cec17e_), .port_680d32a7_(bus_13df4b68_), .port_7e2c6053_(bus_4686658d_), 
  .port_19d5fffb_(Out1_RDY), .port_4ca5ab5a_(repeatRowExpanded_done), .port_6f73ff2c_(consumeRow_done), 
  .port_6a17f116_(reset_done), .port_3c6ad029_(In1_SEND), .DONE(resized_LH2_xy_scheduler_instance_DONE), 
  .RESULT(scheduler), .RESULT_u2119(scheduler_u299), .RESULT_u2120(scheduler_u300), 
  .RESULT_u2121(scheduler_u301), .RESULT_u2122(scheduler_u302), .RESULT_u2123(scheduler_u303), 
  .RESULT_u2124(scheduler_u304), .RESULT_u2125(scheduler_u305), .RESULT_u2126(scheduler_u306), 
  .RESULT_u2127(scheduler_u307), .RESULT_u2128(scheduler_u308), .RESULT_u2129(scheduler_u309), 
  .RESULT_u2130(scheduler_u310), .RESULT_u2131(scheduler_u311), .RESULT_u2132(scheduler_u312), 
  .RESULT_u2133(scheduler_u313), .RESULT_u2134(scheduler_u314), .RESULT_u2135(scheduler_u315), 
  .RESULT_u2136(scheduler_u316));
resized_LH2_xy_stateVar_rowRepeated resized_LH2_xy_stateVar_rowRepeated_1(.bus_2fffcdc9_(CLK), 
  .bus_1df4e7c6_(bus_112f0657_), .bus_543e42b8_(repeatRowExpanded), .bus_3f0e41dd_(repeatRowExpanded_u32), 
  .bus_558d89ec_(reset), .bus_6faa67c2_(16'h1), .bus_45cec17e_(bus_45cec17e_));
resized_LH2_xy_structuralmemory_10a0b0c5_ resized_LH2_xy_structuralmemory_10a0b0c5__1(.CLK_u20(CLK), 
  .bus_5a27453b_(bus_112f0657_), .bus_2abe7aae_(bus_706839bc_), .bus_3da3e1e4_(3'h1), 
  .bus_0a872caa_(bus_1307238a_), .bus_4328a1e0_(bus_0e8f38dd_), .bus_12b5a8c1_(bus_01a9e6ce_), 
  .bus_2b80c1a2_(bus_2b80c1a2_), .bus_2bfcb357_(bus_2bfcb357_));
resized_LH2_xy_reset resized_LH2_xy_reset_instance(.CLK(CLK), .RESET(bus_112f0657_), 
  .GO(reset_go), .DONE(resized_LH2_xy_reset_instance_DONE), .RESULT(reset), .RESULT_u2137(reset_u12), 
  .RESULT_u2138(reset_u13), .RESULT_u2139(reset_u14));
assign bus_7aafd725_=resized_LH2_xy_repeatRowExpanded_instance_DONE&{1{resized_LH2_xy_repeatRowExpanded_instance_DONE}};
resized_LH2_xy_globalreset_physical_0b41fdb2_ resized_LH2_xy_globalreset_physical_0b41fdb2__1(.bus_0a890099_(CLK), 
  .bus_132690ba_(RESET), .bus_112f0657_(bus_112f0657_));
resized_LH2_xy_consumeRow resized_LH2_xy_consumeRow_instance(.CLK(CLK), .RESET(bus_112f0657_), 
  .GO(consumeRow_go), .port_174a8800_(bus_703c1161_), .port_29086a48_(bus_1bceed37_), 
  .port_19cd6551_(bus_4687e307_), .port_21dccef2_(In1_DATA), .DONE(resized_LH2_xy_consumeRow_instance_DONE), 
  .RESULT(consumeRow), .RESULT_u2140(consumeRow_u40), .RESULT_u2145(consumeRow_u41), 
  .RESULT_u2146(consumeRow_u42), .RESULT_u2147(consumeRow_u43), .RESULT_u2148(consumeRow_u44), 
  .RESULT_u2141(consumeRow_u45), .RESULT_u2142(consumeRow_u46), .RESULT_u2143(consumeRow_u47), 
  .RESULT_u2144(consumeRow_u48), .RESULT_u2149(consumeRow_u49));
resized_LH2_xy_stateVar_fsmState_resized_LH2_xy resized_LH2_xy_stateVar_fsmState_resized_LH2_xy_1(.bus_5fb95275_(CLK), 
  .bus_4d57ece6_(bus_112f0657_), .bus_215b8d1b_(scheduler_u300), .bus_46a6a319_(scheduler_u301), 
  .bus_2a450b51_(bus_2a450b51_));
resized_LH2_xy_structuralmemory_57a3ce5d_ resized_LH2_xy_structuralmemory_57a3ce5d__1(.CLK_u21(CLK), 
  .bus_0916e569_(bus_112f0657_), .bus_680f5707_(bus_05401935_), .bus_21a49687_(3'h1), 
  .bus_0aab59c9_(bus_04f85a99_), .bus_3650d95d_(bus_736af7eb_), .bus_1e93c313_(bus_180d93a2_), 
  .bus_0f871660_(bus_0f871660_), .bus_55b75661_(bus_55b75661_));
resized_LH2_xy_stateVar_Out1PortEnable resized_LH2_xy_stateVar_Out1PortEnable_1(.bus_08bf0a8c_(CLK), 
  .bus_5fdb8633_(bus_112f0657_), .bus_0abc9c50_(scheduler_u306), .bus_79cef798_(scheduler_u307), 
  .bus_52d26b67_(bus_52d26b67_));
resized_LH2_xy_simplememoryreferee_7c0f4a30_ resized_LH2_xy_simplememoryreferee_7c0f4a30__1(.bus_10a19532_(CLK), 
  .bus_5397d7e3_(bus_112f0657_), .bus_020ff5a4_(bus_55b75661_), .bus_06009997_(bus_0f871660_), 
  .bus_7a5e2484_(consumeRow_u45), .bus_60ad4ce1_(consumeRow_u47), .bus_0309c2e0_(consumeRow_u46), 
  .bus_0b593446_(3'h1), .bus_05ee34dd_(repeatRowExpanded_u33), .bus_56490b57_(repeatRowExpanded_u35), 
  .bus_5b40276e_(repeatRowExpanded_u34), .bus_7aff8d40_(3'h1), .bus_19414a38_(scheduler_u308), 
  .bus_54364352_(scheduler_u309), .bus_7a0b085e_(3'h1), .bus_180d93a2_(bus_180d93a2_), 
  .bus_05401935_(bus_05401935_), .bus_736af7eb_(bus_736af7eb_), .bus_04f85a99_(bus_04f85a99_), 
  .bus_50563d51_(bus_50563d51_), .bus_4687e307_(bus_4687e307_), .bus_307decb9_(bus_307decb9_), 
  .bus_4686658d_(bus_4686658d_), .bus_13df4b68_(bus_13df4b68_));
endmodule



module resized_LH2_xy_Kicker_45(CLK, RESET, bus_4a33a20e_);
input		CLK;
input		RESET;
output		bus_4a33a20e_;
wire		bus_2713ce3e_;
wire		bus_479a248d_;
reg		kicker_1=1'h0;
reg		kicker_res=1'h0;
wire		bus_7ed5a694_;
reg		kicker_2=1'h0;
wire		bus_1cbbcc2c_;
assign bus_2713ce3e_=~kicker_2;
assign bus_479a248d_=kicker_1&bus_1cbbcc2c_&bus_2713ce3e_;
always @(posedge CLK)
begin
kicker_1<=bus_1cbbcc2c_;
end
always @(posedge CLK)
begin
kicker_res<=bus_479a248d_;
end
assign bus_7ed5a694_=bus_1cbbcc2c_&kicker_1;
always @(posedge CLK)
begin
kicker_2<=bus_7ed5a694_;
end
assign bus_1cbbcc2c_=~RESET;
assign bus_4a33a20e_=kicker_res;
endmodule



module resized_LH2_xy_endianswapper_7a3a6c0f_(endianswapper_7a3a6c0f_in, endianswapper_7a3a6c0f_out);
input	[15:0]	endianswapper_7a3a6c0f_in;
output	[15:0]	endianswapper_7a3a6c0f_out;
assign endianswapper_7a3a6c0f_out=endianswapper_7a3a6c0f_in;
endmodule



module resized_LH2_xy_endianswapper_0dc940a1_(endianswapper_0dc940a1_in, endianswapper_0dc940a1_out);
input	[15:0]	endianswapper_0dc940a1_in;
output	[15:0]	endianswapper_0dc940a1_out;
assign endianswapper_0dc940a1_out=endianswapper_0dc940a1_in;
endmodule



module resized_LH2_xy_stateVar_x(bus_49987487_, bus_5d8644af_, bus_551d1965_, bus_30e7f77b_, bus_75dc4e7a_, bus_7e3885be_, bus_703c1161_);
input		bus_49987487_;
input		bus_5d8644af_;
input		bus_551d1965_;
input	[15:0]	bus_30e7f77b_;
input		bus_75dc4e7a_;
input	[15:0]	bus_7e3885be_;
output	[15:0]	bus_703c1161_;
wire	[15:0]	mux_05ab2089_u0;
reg	[15:0]	stateVar_x_u4=16'h0;
wire	[15:0]	endianswapper_7a3a6c0f_out;
wire	[15:0]	endianswapper_0dc940a1_out;
wire		or_661ebcc7_u0;
assign mux_05ab2089_u0=(bus_551d1965_)?bus_30e7f77b_:16'h0;
always @(posedge bus_49987487_ or posedge bus_5d8644af_)
begin
if (bus_5d8644af_)
stateVar_x_u4<=16'h0;
else if (or_661ebcc7_u0)
stateVar_x_u4<=endianswapper_7a3a6c0f_out;
end
resized_LH2_xy_endianswapper_7a3a6c0f_ resized_LH2_xy_endianswapper_7a3a6c0f__1(.endianswapper_7a3a6c0f_in(mux_05ab2089_u0), 
  .endianswapper_7a3a6c0f_out(endianswapper_7a3a6c0f_out));
assign bus_703c1161_=endianswapper_0dc940a1_out;
resized_LH2_xy_endianswapper_0dc940a1_ resized_LH2_xy_endianswapper_0dc940a1__1(.endianswapper_0dc940a1_in(stateVar_x_u4), 
  .endianswapper_0dc940a1_out(endianswapper_0dc940a1_out));
assign or_661ebcc7_u0=bus_551d1965_|bus_75dc4e7a_;
endmodule



module resized_LH2_xy_endianswapper_232d567d_(endianswapper_232d567d_in, endianswapper_232d567d_out);
input	[31:0]	endianswapper_232d567d_in;
output	[31:0]	endianswapper_232d567d_out;
assign endianswapper_232d567d_out=32'h0;
endmodule



module resized_LH2_xy_endianswapper_3f2f08e7_(endianswapper_3f2f08e7_in, endianswapper_3f2f08e7_out);
input	[31:0]	endianswapper_3f2f08e7_in;
output	[31:0]	endianswapper_3f2f08e7_out;
assign endianswapper_3f2f08e7_out=32'h0;
endmodule



module resized_LH2_xy_stateVar_fsmOldState_resized_LH2_xy(bus_38a242af_, bus_3a6e3652_, bus_54189c3e_, bus_35927e1c_, bus_5bffa9c0_);
input		bus_38a242af_;
input		bus_3a6e3652_;
input		bus_54189c3e_;
input	[31:0]	bus_35927e1c_;
output	[31:0]	bus_5bffa9c0_;
wire	[31:0]	endianswapper_232d567d_out;
wire	[31:0]	endianswapper_3f2f08e7_out;
resized_LH2_xy_endianswapper_232d567d_ resized_LH2_xy_endianswapper_232d567d__1(.endianswapper_232d567d_in(32'h0), 
  .endianswapper_232d567d_out(endianswapper_232d567d_out));
assign bus_5bffa9c0_=32'h0;
resized_LH2_xy_endianswapper_3f2f08e7_ resized_LH2_xy_endianswapper_3f2f08e7__1(.endianswapper_3f2f08e7_in(32'h0), 
  .endianswapper_3f2f08e7_out(endianswapper_3f2f08e7_out));
endmodule



module resized_LH2_xy_endianswapper_60ca2d2f_(endianswapper_60ca2d2f_in, endianswapper_60ca2d2f_out);
input	[31:0]	endianswapper_60ca2d2f_in;
output	[31:0]	endianswapper_60ca2d2f_out;
assign endianswapper_60ca2d2f_out=endianswapper_60ca2d2f_in;
endmodule



module resized_LH2_xy_endianswapper_77b2dcc5_(endianswapper_77b2dcc5_in, endianswapper_77b2dcc5_out);
input	[31:0]	endianswapper_77b2dcc5_in;
output	[31:0]	endianswapper_77b2dcc5_out;
assign endianswapper_77b2dcc5_out=endianswapper_77b2dcc5_in;
endmodule



module resized_LH2_xy_stateVar_Out1MaxTokenIndex(bus_7d661b62_, bus_26c83530_, bus_691cf5a3_, bus_43ea8ee1_, bus_7281aa61_);
input		bus_7d661b62_;
input		bus_26c83530_;
input		bus_691cf5a3_;
input	[31:0]	bus_43ea8ee1_;
output	[31:0]	bus_7281aa61_;
reg	[31:0]	stateVar_Out1MaxTokenIndex_u4=32'h0;
wire	[31:0]	endianswapper_60ca2d2f_out;
wire	[31:0]	endianswapper_77b2dcc5_out;
always @(posedge bus_7d661b62_ or posedge bus_26c83530_)
begin
if (bus_26c83530_)
stateVar_Out1MaxTokenIndex_u4<=32'h0;
else if (bus_691cf5a3_)
stateVar_Out1MaxTokenIndex_u4<=endianswapper_60ca2d2f_out;
end
resized_LH2_xy_endianswapper_60ca2d2f_ resized_LH2_xy_endianswapper_60ca2d2f__1(.endianswapper_60ca2d2f_in(bus_43ea8ee1_), 
  .endianswapper_60ca2d2f_out(endianswapper_60ca2d2f_out));
assign bus_7281aa61_=endianswapper_77b2dcc5_out;
resized_LH2_xy_endianswapper_77b2dcc5_ resized_LH2_xy_endianswapper_77b2dcc5__1(.endianswapper_77b2dcc5_in(stateVar_Out1MaxTokenIndex_u4), 
  .endianswapper_77b2dcc5_out(endianswapper_77b2dcc5_out));
endmodule



module resized_LH2_xy_endianswapper_588803da_(endianswapper_588803da_in, endianswapper_588803da_out);
input	[31:0]	endianswapper_588803da_in;
output	[31:0]	endianswapper_588803da_out;
assign endianswapper_588803da_out=endianswapper_588803da_in;
endmodule



module resized_LH2_xy_endianswapper_24f5942c_(endianswapper_24f5942c_in, endianswapper_24f5942c_out);
input	[31:0]	endianswapper_24f5942c_in;
output	[31:0]	endianswapper_24f5942c_out;
assign endianswapper_24f5942c_out=endianswapper_24f5942c_in;
endmodule



module resized_LH2_xy_stateVar_Out1TokenIndex(bus_71cf89b8_, bus_1502dffb_, bus_2791719c_, bus_29e05130_, bus_3b01d7ce_);
input		bus_71cf89b8_;
input		bus_1502dffb_;
input		bus_2791719c_;
input	[31:0]	bus_29e05130_;
output	[31:0]	bus_3b01d7ce_;
wire	[31:0]	endianswapper_588803da_out;
reg	[31:0]	stateVar_Out1TokenIndex_u4=32'h0;
wire	[31:0]	endianswapper_24f5942c_out;
resized_LH2_xy_endianswapper_588803da_ resized_LH2_xy_endianswapper_588803da__1(.endianswapper_588803da_in(bus_29e05130_), 
  .endianswapper_588803da_out(endianswapper_588803da_out));
assign bus_3b01d7ce_=endianswapper_24f5942c_out;
always @(posedge bus_71cf89b8_ or posedge bus_1502dffb_)
begin
if (bus_1502dffb_)
stateVar_Out1TokenIndex_u4<=32'h0;
else if (bus_2791719c_)
stateVar_Out1TokenIndex_u4<=endianswapper_588803da_out;
end
resized_LH2_xy_endianswapper_24f5942c_ resized_LH2_xy_endianswapper_24f5942c__1(.endianswapper_24f5942c_in(stateVar_Out1TokenIndex_u4), 
  .endianswapper_24f5942c_out(endianswapper_24f5942c_out));
endmodule



module resized_LH2_xy_repeatRowExpanded(CLK, RESET, GO, port_5bf0021c_, port_2dd6a8c5_, port_3f45710a_, port_047547ec_, RESULT, RESULT_u2111, RESULT_u2112, RESULT_u2113, RESULT_u2114, RESULT_u2115, RESULT_u2116, RESULT_u2117, RESULT_u2118, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_5bf0021c_;
input		port_2dd6a8c5_;
input		port_3f45710a_;
input	[15:0]	port_047547ec_;
output		RESULT;
output	[15:0]	RESULT_u2111;
output		RESULT_u2112;
output	[31:0]	RESULT_u2113;
output	[15:0]	RESULT_u2114;
output	[2:0]	RESULT_u2115;
output		RESULT_u2116;
output	[31:0]	RESULT_u2117;
output	[2:0]	RESULT_u2118;
output		DONE;
wire	[15:0]	add;
wire		and_u3596_u0;
reg		and_delayed_u238=1'h0;
wire	[31:0]	add_u473;
wire		and_u3597_u0;
wire	[31:0]	add_u474;
wire		or_u1103_u0;
wire		and_u3598_u0;
reg		reg_51a7597d_u0=1'h0;
wire	[31:0]	add_u475;
reg	[31:0]	syncEnable_u687=32'h0;
wire		lessThan;
wire signed	[31:0]	lessThan_a_signed;
wire signed	[31:0]	lessThan_b_signed;
wire		not_u585_u0;
wire		and_u3599_u0;
wire		and_u3600_u0;
wire		and_u3601_u0;
wire	[31:0]	mux_u359;
wire		or_u1104_u0;
reg		reg_160735b5_u0=1'h0;
assign add=port_5bf0021c_+16'h1;
assign and_u3596_u0=and_u3599_u0&or_u1104_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u238<=1'h0;
else and_delayed_u238<=and_u3596_u0;
end
assign add_u473=mux_u359+32'h0;
assign and_u3597_u0=and_u3596_u0&port_3f45710a_;
assign add_u474=mux_u359+32'h0;
assign or_u1103_u0=and_u3598_u0|RESET;
assign and_u3598_u0=reg_51a7597d_u0&port_2dd6a8c5_;
always @(posedge CLK or posedge and_u3596_u0 or posedge or_u1103_u0)
begin
if (or_u1103_u0)
reg_51a7597d_u0<=1'h0;
else if (and_u3596_u0)
reg_51a7597d_u0<=1'h1;
else reg_51a7597d_u0<=reg_51a7597d_u0;
end
assign add_u475=mux_u359+32'h1;
always @(posedge CLK)
begin
if (and_u3596_u0)
syncEnable_u687<=add_u475;
end
assign lessThan_a_signed=mux_u359;
assign lessThan_b_signed=32'h200;
assign lessThan=lessThan_a_signed<lessThan_b_signed;
assign not_u585_u0=~lessThan;
assign and_u3599_u0=or_u1104_u0&lessThan;
assign and_u3600_u0=or_u1104_u0&not_u585_u0;
assign and_u3601_u0=and_u3600_u0&or_u1104_u0;
assign mux_u359=(reg_160735b5_u0)?32'h0:syncEnable_u687;
assign or_u1104_u0=reg_160735b5_u0|and_delayed_u238;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_160735b5_u0<=1'h0;
else reg_160735b5_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u2111=add;
assign RESULT_u2112=and_u3596_u0;
assign RESULT_u2113=add_u474;
assign RESULT_u2114=port_047547ec_;
assign RESULT_u2115=3'h1;
assign RESULT_u2116=and_u3596_u0;
assign RESULT_u2117=add_u473;
assign RESULT_u2118=3'h1;
assign DONE=and_u3601_u0;
endmodule



module resized_LH2_xy_simplememoryreferee_53c3fe95_(bus_329d11ec_, bus_6055eb84_, bus_23b69ded_, bus_0d07a037_, bus_42291ec9_, bus_4d695e2f_, bus_6f653eab_, bus_7bc2b5e6_, bus_277138ad_, bus_278380fd_, bus_34fe08d6_, bus_01a9e6ce_, bus_706839bc_, bus_0e8f38dd_, bus_1307238a_, bus_551a77e4_, bus_1bceed37_, bus_4bbace21_, bus_768c4387_);
input		bus_329d11ec_;
input		bus_6055eb84_;
input		bus_23b69ded_;
input	[15:0]	bus_0d07a037_;
input		bus_42291ec9_;
input	[15:0]	bus_4d695e2f_;
input	[31:0]	bus_6f653eab_;
input	[2:0]	bus_7bc2b5e6_;
input		bus_277138ad_;
input	[31:0]	bus_278380fd_;
input	[2:0]	bus_34fe08d6_;
output	[15:0]	bus_01a9e6ce_;
output	[31:0]	bus_706839bc_;
output		bus_0e8f38dd_;
output		bus_1307238a_;
output	[2:0]	bus_551a77e4_;
output		bus_1bceed37_;
output	[15:0]	bus_4bbace21_;
output		bus_768c4387_;
wire		and_48326f73_u0;
wire		or_209f369b_u0;
wire		and_48c66f62_u0;
wire		or_2b26a103_u0;
wire		or_5f9c9e39_u0;
wire		not_30e0b2e7_u0;
wire	[15:0]	mux_5b3f6b56_u0;
wire		not_37e52691_u0;
wire	[31:0]	mux_0ee26f39_u0;
reg		done_qual_u195=1'h0;
reg		done_qual_u196_u0=1'h0;
assign and_48326f73_u0=or_209f369b_u0&bus_23b69ded_;
assign or_209f369b_u0=bus_42291ec9_|done_qual_u195;
assign and_48c66f62_u0=or_5f9c9e39_u0&bus_23b69ded_;
assign or_2b26a103_u0=bus_42291ec9_|bus_277138ad_;
assign or_5f9c9e39_u0=bus_277138ad_|done_qual_u196_u0;
assign not_30e0b2e7_u0=~bus_23b69ded_;
assign mux_5b3f6b56_u0=({16{bus_42291ec9_}}&bus_4d695e2f_);
assign not_37e52691_u0=~bus_23b69ded_;
assign bus_01a9e6ce_=mux_5b3f6b56_u0;
assign bus_706839bc_=mux_0ee26f39_u0;
assign bus_0e8f38dd_=bus_42291ec9_;
assign bus_1307238a_=or_2b26a103_u0;
assign bus_551a77e4_=3'h1;
assign bus_1bceed37_=and_48326f73_u0;
assign bus_4bbace21_=bus_0d07a037_;
assign bus_768c4387_=and_48c66f62_u0;
assign mux_0ee26f39_u0=(bus_42291ec9_)?bus_6f653eab_:bus_278380fd_;
always @(posedge bus_329d11ec_)
begin
if (bus_6055eb84_)
done_qual_u195<=1'h0;
else done_qual_u195<=bus_42291ec9_;
end
always @(posedge bus_329d11ec_)
begin
if (bus_6055eb84_)
done_qual_u196_u0<=1'h0;
else done_qual_u196_u0<=bus_277138ad_;
end
endmodule



module resized_LH2_xy_scheduler(CLK, RESET, GO, port_3b0b1e1a_, port_5b3d11e3_, port_5aad7090_, port_598dd3c9_, port_02986e5e_, port_177051de_, port_386b1b7a_, port_680d32a7_, port_7e2c6053_, port_19d5fffb_, port_4ca5ab5a_, port_6f73ff2c_, port_6a17f116_, port_3c6ad029_, RESULT, RESULT_u2119, RESULT_u2120, RESULT_u2121, RESULT_u2122, RESULT_u2123, RESULT_u2124, RESULT_u2125, RESULT_u2126, RESULT_u2127, RESULT_u2128, RESULT_u2129, RESULT_u2130, RESULT_u2131, RESULT_u2132, RESULT_u2133, RESULT_u2134, RESULT_u2135, RESULT_u2136, DONE);
input		CLK;
input		RESET;
input		GO;
input	[31:0]	port_3b0b1e1a_;
input		port_5b3d11e3_;
input	[31:0]	port_5aad7090_;
input	[31:0]	port_598dd3c9_;
input		port_02986e5e_;
input	[15:0]	port_177051de_;
input	[15:0]	port_386b1b7a_;
input		port_680d32a7_;
input	[15:0]	port_7e2c6053_;
input		port_19d5fffb_;
input		port_4ca5ab5a_;
input		port_6f73ff2c_;
input		port_6a17f116_;
input		port_3c6ad029_;
output		RESULT;
output	[31:0]	RESULT_u2119;
output		RESULT_u2120;
output		RESULT_u2121;
output		RESULT_u2122;
output	[31:0]	RESULT_u2123;
output		RESULT_u2124;
output	[31:0]	RESULT_u2125;
output		RESULT_u2126;
output		RESULT_u2127;
output		RESULT_u2128;
output	[31:0]	RESULT_u2129;
output	[2:0]	RESULT_u2130;
output		RESULT_u2131;
output	[15:0]	RESULT_u2132;
output		RESULT_u2133;
output		RESULT_u2134;
output		RESULT_u2135;
output	[15:0]	RESULT_u2136;
output		DONE;
wire	[15:0]	lessThan_a_unsigned;
wire		lessThan;
wire	[15:0]	lessThan_b_unsigned;
wire	[15:0]	equals_a_unsigned;
wire		equals;
wire	[15:0]	equals_b_unsigned;
wire	[15:0]	lessThan_u86_b_unsigned;
wire	[15:0]	lessThan_u86_a_unsigned;
wire		lessThan_u86;
wire		andOp;
wire	[15:0]	equals_u188_b_unsigned;
wire	[15:0]	equals_u188_a_unsigned;
wire		equals_u188;
wire signed	[31:0]	equals_u189_b_signed;
wire		equals_u189;
wire signed	[31:0]	equals_u189_a_signed;
wire		not_u586_u0;
wire		and_u3602_u0;
wire		and_u3603_u0;
wire		andOp_u193;
wire		not_u587_u0;
wire		and_u3604_u0;
wire		and_u3605_u0;
wire		simplePinWrite;
wire		not_u588_u0;
wire		and_u3606_u0;
wire		and_u3607_u0;
wire		simplePinWrite_u516;
wire		and_u3608_u0;
wire		and_u3609_u0;
wire		not_u589_u0;
wire		simplePinWrite_u517;
wire		and_u3610_u0;
reg		reg_351e991f_u0=1'h0;
reg		reg_74967c94_u0=1'h0;
reg		reg_74967c94_result_delayed_u0=1'h0;
reg		reg_3b9cf399_u0=1'h0;
wire		or_u1105_u0;
reg		reg_57b957bf_u0=1'h0;
reg		reg_2c204028_u0=1'h0;
reg		reg_3471a47b_u0=1'h0;
reg		reg_7b991f92_u0=1'h0;
reg		reg_697bf970_u0=1'h0;
reg		reg_3912a11e_u0=1'h0;
reg		reg_5cd550db_u0=1'h0;
reg		reg_51926d82_u0=1'h0;
reg		reg_46946686_u0=1'h0;
reg		reg_29f9ddea_u0=1'h0;
reg		reg_69b415a1_u0=1'h0;
reg		reg_7d7ca566_u0=1'h0;
reg		reg_737da366_u0=1'h0;
reg		reg_5e49b654_u0=1'h0;
reg		reg_1b5b6b45_u0=1'h0;
reg		reg_619c0582_u0=1'h0;
reg		reg_1bf28bed_u0=1'h0;
reg		reg_1b5b6b45_result_delayed_u0=1'h0;
reg		reg_1dc331e7_u0=1'h0;
reg		reg_718f51a9_u0=1'h0;
reg		reg_1b10bf37_u0=1'h0;
reg		reg_44949cbe_u0=1'h0;
reg		reg_3c729058_u0=1'h0;
reg		reg_69b415a1_result_delayed_u0=1'h0;
reg		reg_41edcddd_u0=1'h0;
reg		reg_4ef81ecb_u0=1'h0;
reg		reg_55610952_u0=1'h0;
reg		reg_29f9ddea_result_delayed_u0=1'h0;
reg		reg_787cb445_u0=1'h0;
reg		reg_5d8aa5b1_u0=1'h0;
reg		reg_632eeb10_u0=1'h0;
reg		reg_3736a309_u0=1'h0;
reg		reg_62a002e4_u0=1'h0;
reg		reg_3126cd62_u0=1'h0;
reg		reg_5d242960_u0=1'h0;
reg		reg_4b05af4d_u0=1'h0;
reg		reg_586b6c26_u0=1'h0;
reg		reg_3fddb792_u0=1'h0;
reg		reg_41edcddd_result_delayed_u0=1'h0;
reg		reg_2ddf258d_u0=1'h0;
reg		reg_1af85aaa_u0=1'h0;
reg		reg_09f461a1_u0=1'h0;
reg		reg_25cb699d_u0=1'h0;
reg		reg_1f76a321_u0=1'h0;
reg		reg_6768af3f_u0=1'h0;
reg		reg_2c47481f_u0=1'h0;
reg		reg_04a958f3_u0=1'h0;
reg		reg_7b1fd745_u0=1'h0;
reg		reg_0ac26e9c_u0=1'h0;
reg		reg_1febb7b4_u0=1'h0;
reg		reg_47f4e3ab_u0=1'h0;
reg		reg_1ed112b0_u0=1'h0;
reg		reg_7624ba47_u0=1'h0;
reg		reg_47e56b81_u0=1'h0;
reg		reg_2c204028_result_delayed_u0=1'h0;
reg		reg_3765130d_u0=1'h0;
reg		reg_47c77fae_u0=1'h0;
reg		reg_1dbaf9d0_u0=1'h0;
reg		reg_79ff2594_u0=1'h0;
reg		reg_549798fc_u0=1'h0;
reg		reg_7834905a_u0=1'h0;
reg		reg_408e14fc_u0=1'h0;
reg		reg_7a2b825f_u0=1'h0;
reg		reg_67de13aa_u0=1'h0;
reg		reg_45535925_u0=1'h0;
reg		reg_28e2989b_u0=1'h0;
reg		reg_633a5b40_u0=1'h0;
reg		reg_3471a47b_result_delayed_u0=1'h0;
reg		reg_3912a11e_result_delayed_u0=1'h0;
reg		reg_7a5ce622_u0=1'h0;
reg		reg_5b32ffb2_u0=1'h0;
reg		reg_71b3a931_u0=1'h0;
reg		reg_23c90b4d_u0=1'h0;
reg		reg_19b1e534_u0=1'h0;
reg		reg_18b39c34_u0=1'h0;
reg		reg_0ac6524e_u0=1'h0;
reg		reg_4a991a10_u0=1'h0;
reg		reg_2bd5f75e_u0=1'h0;
reg		reg_005750dc_u0=1'h0;
reg		reg_67de13aa_result_delayed_u0=1'h0;
reg		reg_029c8613_u0=1'h0;
reg		reg_039f5f0f_u0=1'h0;
reg		reg_31ec057e_u0=1'h0;
reg		reg_1742dbd1_u0=1'h0;
reg		reg_28e17c75_u0=1'h0;
reg		reg_7fe56773_u0=1'h0;
reg		reg_7dcd9154_u0=1'h0;
reg		reg_15d1894b_u0=1'h0;
reg		reg_66fd0261_u0=1'h0;
reg		reg_25cb699d_result_delayed_u0=1'h0;
reg		reg_408e14fc_result_delayed_u0=1'h0;
reg		reg_1dbaf9d0_result_delayed_u0=1'h0;
reg		reg_34478ce7_u0=1'h0;
reg		reg_7b86d327_u0=1'h0;
reg		reg_44949cbe_result_delayed_u0=1'h0;
reg		reg_446bb0cd_u0=1'h0;
reg		reg_449ea438_u0=1'h0;
reg		reg_32d59a7c_u0=1'h0;
reg		reg_5fce0764_u0=1'h0;
reg		reg_7432b099_u0=1'h0;
reg		reg_3471a47b_result_delayed_result_delayed_u0=1'h0;
reg		reg_3de6494b_u0=1'h0;
reg		reg_527dd6cc_u0=1'h0;
reg		reg_6fd8576b_u0=1'h0;
reg		reg_392f0d9b_u0=1'h0;
reg		reg_4a825e39_u0=1'h0;
reg		reg_2c204028_result_delayed_result_delayed_u0=1'h0;
reg		reg_4da6e166_u0=1'h0;
reg		reg_713e21fb_u0=1'h0;
reg		reg_5d8aa5b1_result_delayed_u0=1'h0;
reg		reg_42c05205_u0=1'h0;
reg		reg_449ea438_result_delayed_u0=1'h0;
reg		reg_11f3093e_u0=1'h0;
reg		reg_4c2ecce3_u0=1'h0;
reg		reg_350541ca_u0=1'h0;
reg		reg_7cb11462_u0=1'h0;
reg		reg_45a71573_u0=1'h0;
reg		reg_28bd586b_u0=1'h0;
reg		reg_44949cbe_result_delayed_result_delayed_u0=1'h0;
reg		reg_368fce58_u0=1'h0;
reg		reg_039aa343_u0=1'h0;
reg		reg_4c87c45c_u0=1'h0;
reg		reg_062cdef7_u0=1'h0;
reg		reg_3a1feec1_u0=1'h0;
reg		reg_6f802f62_u0=1'h0;
reg		reg_73ced32a_u0=1'h0;
reg		reg_1cc24c27_u0=1'h0;
reg		reg_7b9f9b79_u0=1'h0;
reg		reg_2ae45e03_u0=1'h0;
reg		reg_1b2287cc_u0=1'h0;
reg		reg_3d4fe5be_u0=1'h0;
reg		reg_3afa1e08_u0=1'h0;
reg		reg_1ba0d353_u0=1'h0;
reg		reg_1b78238d_u0=1'h0;
reg		reg_2632face_u0=1'h0;
reg		reg_7fca9f36_u0=1'h0;
reg		reg_7dd95126_u0=1'h0;
reg		reg_0993b092_u0=1'h0;
reg		reg_12299b2b_u0=1'h0;
reg		reg_7ce161e2_u0=1'h0;
reg		reg_7ce161e2_result_delayed_u0=1'h0;
reg		reg_3a62176b_u0=1'h0;
reg		reg_029c8613_result_delayed_u0=1'h0;
reg		reg_01539059_u0=1'h0;
reg		reg_4bc316c8_u0=1'h0;
reg		reg_0af8dff3_u0=1'h0;
reg		reg_69ccc0c7_u0=1'h0;
reg		reg_7432b099_result_delayed_u0=1'h0;
reg		reg_3b2ea222_u0=1'h0;
reg		reg_5792329f_u0=1'h0;
reg		reg_46946686_result_delayed_u0=1'h0;
reg		reg_67e61ef6_u0=1'h0;
reg		reg_3471a47b_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_1b5b6b45_result_delayed_result_delayed_u0=1'h0;
reg		reg_70705567_u0=1'h0;
reg		reg_1324a63d_u0=1'h0;
reg		reg_2ae45e03_result_delayed_u0=1'h0;
reg		reg_3afa1e08_result_delayed_u0=1'h0;
reg		reg_71d3e4cd_u0=1'h0;
reg		reg_6e167f08_u0=1'h0;
reg		reg_4012210d_u0=1'h0;
reg		reg_0127d038_u0=1'h0;
reg		reg_30e129c3_u0=1'h0;
reg		reg_2b525e7b_u0=1'h0;
reg		reg_134a2263_u0=1'h0;
reg		reg_70705567_result_delayed_u0=1'h0;
reg		reg_2901482a_u0=1'h0;
reg		reg_0924240b_u0=1'h0;
reg		reg_0188e8a7_u0=1'h0;
reg		reg_3afa1e08_result_delayed_result_delayed_u0=1'h0;
reg		reg_63aaa29e_u0=1'h0;
reg		reg_77462671_u0=1'h0;
reg		reg_408e14fc_result_delayed_result_delayed_u0=1'h0;
reg		reg_446bb0cd_result_delayed_u0=1'h0;
reg		reg_527dd6cc_result_delayed_u0=1'h0;
reg		reg_05b504f5_u0=1'h0;
reg		reg_7b991f92_result_delayed_u0=1'h0;
reg		reg_7fa5f2e1_u0=1'h0;
reg		reg_5fc7b281_u0=1'h0;
reg		reg_08cf2d88_u0=1'h0;
reg		reg_2d083c40_u0=1'h0;
reg		reg_62aecfe4_u0=1'h0;
wire		and_u3611_u0;
reg		reg_449ea438_result_delayed_result_delayed_u0=1'h0;
reg		reg_0525586a_u0=1'h0;
reg		reg_25cb699d_result_delayed_result_delayed_u0=1'h0;
reg		reg_4f8742d5_u0=1'h0;
reg		reg_350541ca_result_delayed_u0=1'h0;
reg		reg_44b53de6_u0=1'h0;
reg		reg_6a945bc0_u0=1'h0;
reg		reg_5d8aa5b1_result_delayed_result_delayed_u0=1'h0;
reg		reg_4b05af4d_result_delayed_u0=1'h0;
reg		reg_619c0582_result_delayed_u0=1'h0;
reg		reg_60f8cda6_u0=1'h0;
reg		reg_1801415e_u0=1'h0;
reg		reg_1ec2c3a2_u0=1'h0;
reg		reg_74967c94_result_delayed_result_delayed_u0=1'h0;
reg		reg_12bc27dd_u0=1'h0;
reg		reg_3d2ae849_u0=1'h0;
reg		reg_7a349f51_u0=1'h0;
reg		reg_62aecfe4_result_delayed_u0=1'h0;
reg		reg_47e56b81_result_delayed_u0=1'h0;
reg		reg_0ac26e9c_result_delayed_u0=1'h0;
reg		reg_2ce4bd89_u0=1'h0;
reg		reg_27d7caa5_u0=1'h0;
reg		reg_6a850ff6_u0=1'h0;
reg		reg_12bc27dd_result_delayed_u0=1'h0;
reg		reg_7f9742e2_u0=1'h0;
reg		reg_719ae8ef_u0=1'h0;
reg		reg_6efe4388_u0=1'h0;
reg		reg_1801415e_result_delayed_u0=1'h0;
reg		reg_1cb40934_u0=1'h0;
reg		reg_351e991f_result_delayed_u0=1'h0;
reg		reg_10d31157_u0=1'h0;
reg		reg_2377f2f2_u0=1'h0;
reg		reg_61ecb46b_u0=1'h0;
reg		reg_602c59ab_u0=1'h0;
reg		reg_41edcddd_result_delayed_result_delayed_u0=1'h0;
reg		reg_54ab7523_u0=1'h0;
reg		reg_385515de_u0=1'h0;
reg		reg_6a945bc0_result_delayed_u0=1'h0;
reg		reg_03b7ae24_u0=1'h0;
reg		reg_3765130d_result_delayed_u0=1'h0;
reg		reg_2b525e7b_result_delayed_u0=1'h0;
reg		reg_7121f4b8_u0=1'h0;
reg		reg_52798be3_u0=1'h0;
reg		reg_5e49b654_result_delayed_u0=1'h0;
reg		reg_2fe53643_u0=1'h0;
reg		reg_2c47481f_result_delayed_u0=1'h0;
reg		reg_37b15a18_u0=1'h0;
reg		reg_6efe4388_result_delayed_u0=1'h0;
reg		reg_3052e1e7_u0=1'h0;
reg		reg_5236af83_u0=1'h0;
reg		reg_7b1fd745_result_delayed_u0=1'h0;
reg		reg_010e94b1_u0=1'h0;
reg		reg_3c844144_u0=1'h0;
reg		reg_0af8dff3_result_delayed_u0=1'h0;
reg		reg_4ff65e34_u0=1'h0;
reg		reg_69b415a1_result_delayed_result_delayed_u0=1'h0;
reg		reg_69f58839_u0=1'h0;
reg		reg_719ae8ef_result_delayed_u0=1'h0;
reg		reg_1ed112b0_result_delayed_u0=1'h0;
reg		reg_16e37f2c_u0=1'h0;
reg		reg_3fddb792_result_delayed_u0=1'h0;
reg		reg_1dca001c_u0=1'h0;
reg		reg_08cf2d88_result_delayed_u0=1'h0;
reg		reg_43dd6207_u0=1'h0;
reg		reg_0bd5de0a_u0=1'h0;
reg		reg_3db3d453_u0=1'h0;
reg		reg_3765130d_result_delayed_result_delayed_u0=1'h0;
reg		reg_713e21fb_result_delayed_u0=1'h0;
reg		reg_1dbaf9d0_result_delayed_result_delayed_u0=1'h0;
reg		reg_13ea2607_u0=1'h0;
reg		reg_0924240b_result_delayed_u0=1'h0;
reg		reg_3c729058_result_delayed_u0=1'h0;
reg		and_delayed_u239=1'h0;
reg		reg_005750dc_result_delayed_u0=1'h0;
reg		reg_568a337f_u0=1'h0;
reg		reg_1742dbd1_result_delayed_u0=1'h0;
reg		reg_26a95b50_u0=1'h0;
reg		reg_2fbb9e45_u0=1'h0;
reg		reg_193758c8_u0=1'h0;
reg		reg_713c4f38_u0=1'h0;
reg		reg_49656763_u0=1'h0;
reg		reg_6bfaddf3_u0=1'h0;
reg		reg_1cc24c27_result_delayed_u0=1'h0;
reg		reg_582b1a27_u0=1'h0;
reg		reg_527dd6cc_result_delayed_result_delayed_u0=1'h0;
reg		reg_787cb445_result_delayed_u0=1'h0;
reg		reg_01539059_result_delayed_u0=1'h0;
reg		reg_622e780a_u0=1'h0;
reg		reg_5cd550db_result_delayed_u0=1'h0;
reg		reg_40f3fed8_u0=1'h0;
reg		reg_2e453868_u0=1'h0;
reg		reg_2d501b7f_u0=1'h0;
reg		reg_449ea438_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_1611b424_u0=1'h0;
reg		reg_0f0fdd38_u0=1'h0;
reg		reg_582b1a27_result_delayed_u0=1'h0;
reg		reg_1b10bf37_result_delayed_u0=1'h0;
reg		reg_6a83a8be_u0=1'h0;
reg		reg_713e21fb_result_delayed_result_delayed_u0=1'h0;
reg		reg_37b15a18_result_delayed_u0=1'h0;
reg		reg_12e4f0a0_u0=1'h0;
reg		reg_29f9ddea_result_delayed_result_delayed_u0=1'h0;
reg		reg_787cb445_result_delayed_result_delayed_u0=1'h0;
reg		reg_50e10aad_u0=1'h0;
reg		reg_0b45c90a_u0=1'h0;
reg		reg_0820ce74_u0=1'h0;
reg		reg_4c4df618_u0=1'h0;
reg		reg_55610952_result_delayed_u0=1'h0;
reg		reg_7b1fd745_result_delayed_result_delayed_u0=1'h0;
reg		reg_79ff2594_result_delayed_u0=1'h0;
reg		reg_1a8ce0d2_u0=1'h0;
reg		reg_190e5b6d_u0=1'h0;
reg		reg_286c1a08_u0=1'h0;
reg		reg_17bf09db_u0=1'h0;
reg		reg_15fe439b_u0=1'h0;
reg		reg_7624ba47_result_delayed_u0=1'h0;
reg		reg_42fabc9d_u0=1'h0;
reg		reg_1130ef58_u0=1'h0;
reg		reg_6a83a8be_result_delayed_u0=1'h0;
reg		reg_47f4e3ab_result_delayed_u0=1'h0;
reg		reg_719347fd_u0=1'h0;
reg		reg_6a945bc0_result_delayed_result_delayed_u0=1'h0;
reg		reg_7a2b825f_result_delayed_u0=1'h0;
reg		reg_049d62ec_u0=1'h0;
reg		reg_1795d1e7_u0=1'h0;
reg		reg_62a002e4_result_delayed_u0=1'h0;
reg		reg_4650dc26_u0=1'h0;
reg		reg_5b32ffb2_result_delayed_u0=1'h0;
reg		reg_1f76a321_result_delayed_u0=1'h0;
reg		reg_2dc36fb8_u0=1'h0;
reg		reg_737be907_u0=1'h0;
reg		reg_09f461a1_result_delayed_u0=1'h0;
reg		reg_65dbefa4_u0=1'h0;
reg		reg_51cd934d_u0=1'h0;
reg		reg_51004f81_u0=1'h0;
reg		reg_69ccc0c7_result_delayed_u0=1'h0;
reg		reg_0924240b_result_delayed_result_delayed_u0=1'h0;
reg		reg_549798fc_result_delayed_u0=1'h0;
reg		reg_67e61ef6_result_delayed_u0=1'h0;
reg		reg_69f58839_result_delayed_u0=1'h0;
reg		reg_3d2ae849_result_delayed_u0=1'h0;
reg		reg_1b5b6b45_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_41edcddd_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_1dbaf9d0_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_6fd8576b_result_delayed_u0=1'h0;
reg		reg_190e5b6d_result_delayed_u0=1'h0;
reg		reg_26a95b50_result_delayed_u0=1'h0;
reg		reg_57b957bf_result_delayed_u0=1'h0;
reg		reg_549798fc_result_delayed_result_delayed_u0=1'h0;
reg		reg_44b53de6_result_delayed_u0=1'h0;
reg		reg_2fe53643_result_delayed_u0=1'h0;
reg		reg_010e94b1_result_delayed_u0=1'h0;
reg		reg_7ce161e2_result_delayed_result_delayed_u0=1'h0;
reg		reg_092d4389_u0=1'h0;
reg		reg_7cb11462_result_delayed_u0=1'h0;
reg		reg_633a799d_u0=1'h0;
reg		reg_2ded6345_u0=1'h0;
reg		reg_0db7cb1d_u0=1'h0;
reg		reg_7fe56773_result_delayed_u0=1'h0;
reg		reg_08ab9607_u0=1'h0;
reg		reg_37d2817c_u0=1'h0;
reg		reg_12247897_u0=1'h0;
reg		reg_4c4df618_result_delayed_u0=1'h0;
reg		reg_67e61ef6_result_delayed_result_delayed_u0=1'h0;
reg		reg_60d46663_u0=1'h0;
reg		reg_2a6d54d5_u0=1'h0;
reg		reg_0f03e5b9_u0=1'h0;
reg		reg_5792329f_result_delayed_u0=1'h0;
reg		reg_2632face_result_delayed_u0=1'h0;
reg		reg_2bd5f75e_result_delayed_u0=1'h0;
reg		reg_617de3bd_u0=1'h0;
reg		reg_26a95b50_result_delayed_result_delayed_u0=1'h0;
reg		reg_6f802f62_result_delayed_u0=1'h0;
reg		reg_15fe439b_result_delayed_u0=1'h0;
reg		reg_0ac6524e_result_delayed_u0=1'h0;
reg		reg_5e962850_u0=1'h0;
reg		reg_4012210d_result_delayed_u0=1'h0;
reg		reg_07488981_u0=1'h0;
reg		reg_4874c2bd_u0=1'h0;
reg		reg_582b1a27_result_delayed_result_delayed_u0=1'h0;
reg		reg_0127d038_result_delayed_u0=1'h0;
reg		reg_3ef9b436_u0=1'h0;
reg		reg_4f8742d5_result_delayed_u0=1'h0;
reg		reg_7121f4b8_result_delayed_u0=1'h0;
reg		reg_27d7caa5_result_delayed_u0=1'h0;
reg		reg_18b39c34_result_delayed_u0=1'h0;
reg		reg_1554b782_u0=1'h0;
reg		reg_2c47481f_result_delayed_result_delayed_u0=1'h0;
reg		reg_1af85aaa_result_delayed_u0=1'h0;
reg		reg_446bb0cd_result_delayed_result_delayed_u0=1'h0;
reg		reg_54ab7523_result_delayed_u0=1'h0;
reg		reg_69e5773a_u0=1'h0;
reg		reg_31ec057e_result_delayed_u0=1'h0;
reg		reg_3471a47b_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_713e21fb_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_072dadc1_u0=1'h0;
reg		reg_17bf09db_result_delayed_u0=1'h0;
reg		reg_70705567_result_delayed_result_delayed_u0=1'h0;
reg		reg_23c90b4d_result_delayed_u0=1'h0;
reg		reg_0224b0d4_u0=1'h0;
reg		reg_3c1b12e8_u0=1'h0;
reg		reg_27d7caa5_result_delayed_result_delayed_u0=1'h0;
reg		reg_408e14fc_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_12247897_result_delayed_u0=1'h0;
reg		reg_486de694_u0=1'h0;
reg		reg_11cd6f36_u0=1'h0;
reg		reg_47f4e3ab_result_delayed_result_delayed_u0=1'h0;
reg		reg_11f3093e_result_delayed_u0=1'h0;
reg		reg_713c4f38_result_delayed_u0=1'h0;
reg		reg_5dc782c5_u0=1'h0;
reg		reg_1b2287cc_result_delayed_u0=1'h0;
reg		reg_1dca001c_result_delayed_u0=1'h0;
reg		reg_46b7b9ba_u0=1'h0;
reg		reg_3de6494b_result_delayed_u0=1'h0;
reg		reg_7f9742e2_result_delayed_u0=1'h0;
reg		reg_6a948183_u0=1'h0;
reg		reg_66fd0261_result_delayed_u0=1'h0;
reg		reg_5fc7b281_result_delayed_u0=1'h0;
reg		reg_134a2263_result_delayed_u0=1'h0;
reg		reg_7a2b825f_result_delayed_result_delayed_u0=1'h0;
reg		reg_36c619e0_u0=1'h0;
reg		reg_719ae8ef_result_delayed_result_delayed_u0=1'h0;
wire		and_u3612_u0;
reg		reg_51926d82_result_delayed_u0=1'h0;
reg		reg_71134e38_u0=1'h0;
reg		reg_7b86d327_result_delayed_u0=1'h0;
reg		reg_28e2989b_result_delayed_u0=1'h0;
reg		reg_11f3093e_result_delayed_result_delayed_u0=1'h0;
reg		reg_0820ce74_result_delayed_u0=1'h0;
reg		reg_1554b782_result_delayed_u0=1'h0;
reg		reg_71d3e4cd_result_delayed_u0=1'h0;
reg		reg_5d242960_result_delayed_u0=1'h0;
reg		reg_50e10aad_result_delayed_u0=1'h0;
reg		reg_7ee659a2_u0=1'h0;
reg		reg_1febb7b4_result_delayed_u0=1'h0;
reg		reg_28e17c75_result_delayed_u0=1'h0;
reg		reg_4fad7ce4_u0=1'h0;
reg		reg_718f51a9_result_delayed_u0=1'h0;
reg		reg_1dc331e7_result_delayed_u0=1'h0;
reg		reg_2fbb9e45_result_delayed_u0=1'h0;
reg		reg_47c77fae_result_delayed_u0=1'h0;
reg		reg_350541ca_result_delayed_result_delayed_u0=1'h0;
reg		reg_1bf28bed_result_delayed_u0=1'h0;
reg		reg_79ff2594_result_delayed_result_delayed_u0=1'h0;
reg		reg_57e6dcb6_u0=1'h0;
reg		reg_63aaa29e_result_delayed_u0=1'h0;
reg		reg_05b504f5_result_delayed_u0=1'h0;
reg		reg_2bd5f75e_result_delayed_result_delayed_u0=1'h0;
reg		reg_51004f81_result_delayed_u0=1'h0;
reg		reg_5d8aa5b1_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_71134e38_result_delayed_u0=1'h0;
reg		reg_385515de_result_delayed_u0=1'h0;
reg		reg_60d46663_result_delayed_u0=1'h0;
reg		reg_62aecfe4_result_delayed_result_delayed_u0=1'h0;
reg		reg_08cf2d88_result_delayed_result_delayed_u0=1'h0;
reg		reg_04a958f3_result_delayed_u0=1'h0;
reg		reg_632eeb10_result_delayed_u0=1'h0;
reg		reg_2ddf258d_result_delayed_u0=1'h0;
reg		reg_549798fc_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_1324a63d_result_delayed_u0=1'h0;
reg		reg_7dd95126_result_delayed_u0=1'h0;
reg		reg_3a62176b_result_delayed_u0=1'h0;
reg		reg_2499b3e8_u0=1'h0;
reg		reg_4f8742d5_result_delayed_result_delayed_u0=1'h0;
reg		reg_15d1894b_result_delayed_u0=1'h0;
reg		reg_47e56b81_result_delayed_result_delayed_u0=1'h0;
reg		reg_30e129c3_result_delayed_u0=1'h0;
reg		reg_46b7b9ba_result_delayed_u0=1'h0;
reg		reg_005750dc_result_delayed_result_delayed_u0=1'h0;
reg		reg_5236af83_result_delayed_u0=1'h0;
reg		reg_029c8613_result_delayed_result_delayed_u0=1'h0;
reg		reg_69b415a1_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_6a850ff6_result_delayed_u0=1'h0;
reg		reg_1f3d20af_u0=1'h0;
reg		reg_4ef81ecb_result_delayed_u0=1'h0;
reg		reg_7a5ce622_result_delayed_u0=1'h0;
reg		reg_6efe4388_result_delayed_result_delayed_u0=1'h0;
reg		reg_7b991f92_result_delayed_result_delayed_u0=1'h0;
reg		reg_12bc27dd_result_delayed_result_delayed_u0=1'h0;
reg		reg_4bc316c8_result_delayed_u0=1'h0;
reg		reg_33a8b808_u0=1'h0;
reg		reg_63cbe06a_u0=1'h0;
reg		reg_1795d1e7_result_delayed_u0=1'h0;
reg		reg_3126cd62_result_delayed_u0=1'h0;
reg		reg_37b15a18_result_delayed_result_delayed_u0=1'h0;
reg		reg_1324a63d_result_delayed_result_delayed_u0=1'h0;
reg		reg_3db3d453_result_delayed_u0=1'h0;
reg		reg_697bf970_result_delayed_u0=1'h0;
reg		reg_51cd934d_result_delayed_u0=1'h0;
reg		reg_1554b782_result_delayed_result_delayed_u0=1'h0;
reg		reg_0f0fdd38_result_delayed_u0=1'h0;
reg		reg_45a71573_result_delayed_u0=1'h0;
reg		reg_12e4f0a0_result_delayed_u0=1'h0;
reg		reg_34478ce7_result_delayed_u0=1'h0;
reg		reg_3b9cf399_result_delayed_u0=1'h0;
reg		reg_1ec2c3a2_result_delayed_u0=1'h0;
reg		reg_4fad7ce4_result_delayed_u0=1'h0;
reg		reg_16e37f2c_result_delayed_u0=1'h0;
reg		reg_25cb699d_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_19b1e534_result_delayed_u0=1'h0;
reg		reg_787cb445_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_6768af3f_result_delayed_u0=1'h0;
reg		reg_7d7ca566_result_delayed_u0=1'h0;
reg		reg_65dbefa4_result_delayed_u0=1'h0;
reg		reg_0924240b_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_40f3fed8_result_delayed_u0=1'h0;
reg		reg_0f03e5b9_result_delayed_u0=1'h0;
reg		reg_7cb11462_result_delayed_result_delayed_u0=1'h0;
reg		reg_29f9ddea_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_2bd5f75e_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_52798be3_result_delayed_u0=1'h0;
reg		reg_09f461a1_result_delayed_result_delayed_u0=1'h0;
reg		reg_633a5b40_result_delayed_u0=1'h0;
reg		reg_1ba0d353_result_delayed_u0=1'h0;
reg		reg_7b9f9b79_result_delayed_u0=1'h0;
reg		reg_10d31157_result_delayed_u0=1'h0;
reg		reg_368fce58_result_delayed_u0=1'h0;
reg		reg_2ae45e03_result_delayed_result_delayed_u0=1'h0;
reg		reg_79ff2594_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_12299b2b_result_delayed_u0=1'h0;
reg		reg_0bd5de0a_result_delayed_u0=1'h0;
reg		reg_32d59a7c_result_delayed_u0=1'h0;
reg		reg_7834905a_result_delayed_u0=1'h0;
reg		reg_039f5f0f_result_delayed_u0=1'h0;
reg		reg_04a958f3_result_delayed_result_delayed_u0=1'h0;
reg		reg_4ef81ecb_result_delayed_result_delayed_u0=1'h0;
wire		or_u1106_u0;
wire		mux_u360;
reg		reg_787cb445_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_1801415e_result_delayed_result_delayed_u0=1'h0;
reg		reg_11cd6f36_result_delayed_u0=1'h0;
wire		mux_u361_u0;
wire		or_u1107_u0;
wire		or_u1108_u0;
wire	[31:0]	mux_u362_u0;
reg		reg_4e481e21_u0=1'h0;
reg		reg_2258ca11_u0=1'h0;
wire		or_u1109_u0;
wire		and_u3613_u0;
wire		or_u1110_u0;
wire		or_u1111_u0;
reg		reg_4e481e21_result_delayed_u0=1'h0;
reg		reg_3a07cc10_u0=1'h0;
wire		or_u1112_u0;
wire		and_u3614_u0;
reg		reg_4e481e21_result_delayed_result_delayed_u0=1'h0;
wire		and_u3615_u0;
reg		and_delayed_u240_u0=1'h0;
wire		or_u1113_u0;
wire		and_u3616_u0;
wire signed	[31:0]	equals_u190_b_signed;
wire		equals_u190;
wire signed	[31:0]	equals_u190_a_signed;
wire		and_u3617_u0;
wire		not_u590_u0;
wire		and_u3618_u0;
wire		and_u3619_u0;
wire		not_u591_u0;
wire		and_u3620_u0;
wire		lessThan_u87;
wire signed	[31:0]	lessThan_u87_a_signed;
wire signed	[31:0]	lessThan_u87_b_signed;
wire		not_u592_u0;
wire		and_u3621_u0;
wire		and_u3622_u0;
wire		and_u3623_u0;
wire		not_u593_u0;
wire		and_u3624_u0;
wire	[31:0]	add;
wire		and_u3625_u0;
wire		simplePinWrite_u518;
wire	[15:0]	simplePinWrite_u519;
wire	[15:0]	simplePinWrite_u520;
wire	[31:0]	add_u476;
reg	[15:0]	syncEnable_u688=16'h0;
wire		and_u3626_u0;
reg		and_delayed_u241_u0=1'h0;
reg		reg_22db32bc_u0=1'h0;
wire		and_u3627_u0;
wire	[15:0]	mux_u363_u0;
reg	[15:0]	syncEnable_u689_u0=16'h0;
wire		and_u3628_u0;
reg		and_delayed_u242_u0=1'h0;
wire	[15:0]	mux_u364_u0;
wire		and_u3629_u0;
reg		and_delayed_u243_u0=1'h0;
wire	[31:0]	mux_u365_u0;
reg	[15:0]	syncEnable_u690_u0=16'h0;
reg	[31:0]	syncEnable_u691_u0=32'h0;
wire	[31:0]	mux_u366_u0;
reg		reg_10a5074b_u0=1'h0;
wire	[15:0]	mux_u367_u0;
reg	[31:0]	syncEnable_u692_u0=32'h0;
wire		and_u3630_u0;
reg		and_delayed_u244_u0=1'h0;
reg	[15:0]	syncEnable_u693_u0=16'h0;
wire		and_u3631_u0;
reg	[15:0]	syncEnable_u694_u0=16'h0;
wire		and_u3632_u0;
reg		and_delayed_u245_u0=1'h0;
wire		and_u3633_u0;
wire	[31:0]	mux_u368_u0;
reg	[31:0]	syncEnable_u695_u0=32'h0;
reg		and_delayed_u246_u0=1'h0;
wire	[15:0]	mux_u369_u0;
wire	[31:0]	mux_u370_u0;
wire		or_u1114_u0;
wire	[31:0]	latch_512b7f83_out;
reg	[31:0]	latch_512b7f83_reg=32'h0;
reg	[15:0]	latch_57dc3c15_reg=16'h0;
wire	[15:0]	latch_57dc3c15_out;
wire		or_u1115_u0;
wire		mux_u371_u0;
reg		block_GO_delayed_u12=1'h0;
wire	[31:0]	mux_u372_u0;
wire		or_u1116_u0;
wire		or_u1117_u0;
wire		mux_u373_u0;
wire		and_u3634_u0;
reg		loopControl_u9=1'h0;
wire		or_u1118_u0;
reg		syncEnable_u696_u0=1'h0;
reg	[15:0]	fbReg_Out1Portvalue_u4=16'h0;
reg	[31:0]	fbReg_temp_fsmOldState_resized_LH2_xy_7_u0=32'h0;
wire	[31:0]	mux_u374_u0;
wire	[15:0]	mux_u375_u0;
wire		or_u1119_u0;
wire		mux_u376_u0;
wire		mux_u377_u0;
wire		or_u1120_u0;
wire		or_u1121_u0;
wire		or_u1122_u0;
wire	[31:0]	mux_u378_u0;
wire	[31:0]	mux_u379_u0;
wire		or_u1123_u0;
reg		reg_7a06e94d_u0=1'h0;
reg		reg_7a06e94d_result_delayed_u0=1'h0;
assign lessThan_a_unsigned=port_177051de_;
assign lessThan_b_unsigned=16'h80;
assign lessThan=lessThan_a_unsigned<lessThan_b_unsigned;
assign equals_a_unsigned=port_177051de_;
assign equals_b_unsigned=16'h80;
assign equals=equals_a_unsigned==equals_b_unsigned;
assign lessThan_u86_a_unsigned=port_386b1b7a_;
assign lessThan_u86_b_unsigned=16'h4;
assign lessThan_u86=lessThan_u86_a_unsigned<lessThan_u86_b_unsigned;
assign andOp=equals&lessThan_u86;
assign equals_u188_a_unsigned=port_386b1b7a_;
assign equals_u188_b_unsigned=16'h4;
assign equals_u188=equals_u188_a_unsigned==equals_u188_b_unsigned;
assign equals_u189_a_signed={31'b0, port_5b3d11e3_};
assign equals_u189_b_signed=32'h0;
assign equals_u189=equals_u189_a_signed==equals_u189_b_signed;
assign not_u586_u0=~equals_u189;
assign and_u3602_u0=and_u3634_u0&equals_u189;
assign and_u3603_u0=and_u3634_u0&not_u586_u0;
assign andOp_u193=lessThan&port_3c6ad029_;
assign not_u587_u0=~andOp_u193;
assign and_u3604_u0=and_u3616_u0&andOp_u193;
assign and_u3605_u0=and_u3616_u0&not_u587_u0;
assign simplePinWrite=and_u3614_u0&{1{and_u3614_u0}};
assign not_u588_u0=~andOp;
assign and_u3606_u0=and_u3613_u0&andOp;
assign and_u3607_u0=and_u3613_u0&not_u588_u0;
assign simplePinWrite_u516=and_u3611_u0&{1{and_u3611_u0}};
assign and_u3608_u0=and_u3612_u0&equals_u188;
assign and_u3609_u0=and_u3612_u0&not_u589_u0;
assign not_u589_u0=~equals_u188;
assign simplePinWrite_u517=and_u3610_u0&{1{and_u3610_u0}};
assign and_u3610_u0=and_u3608_u0&and_u3612_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_351e991f_u0<=1'h0;
else reg_351e991f_u0<=reg_71b3a931_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_74967c94_u0<=1'h0;
else reg_74967c94_u0<=reg_6fd8576b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_74967c94_result_delayed_u0<=1'h0;
else reg_74967c94_result_delayed_u0<=reg_74967c94_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3b9cf399_u0<=1'h0;
else reg_3b9cf399_u0<=reg_0127d038_result_delayed_u0;
end
assign or_u1105_u0=reg_7dcd9154_u0|reg_4c2ecce3_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_57b957bf_u0<=1'h0;
else reg_57b957bf_u0<=reg_7432b099_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2c204028_u0<=1'h0;
else reg_2c204028_u0<=reg_01539059_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3471a47b_u0<=1'h0;
else reg_3471a47b_u0<=reg_1795d1e7_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7b991f92_u0<=1'h0;
else reg_7b991f92_u0<=reg_2bd5f75e_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_697bf970_u0<=1'h0;
else reg_697bf970_u0<=reg_0db7cb1d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3912a11e_u0<=1'h0;
else reg_3912a11e_u0<=reg_6bfaddf3_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5cd550db_u0<=1'h0;
else reg_5cd550db_u0<=reg_03b7ae24_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_51926d82_u0<=1'h0;
else reg_51926d82_u0<=reg_737da366_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_46946686_u0<=1'h0;
else reg_46946686_u0<=reg_5fce0764_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_29f9ddea_u0<=1'h0;
else reg_29f9ddea_u0<=reg_2c204028_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_69b415a1_u0<=1'h0;
else reg_69b415a1_u0<=reg_619c0582_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7d7ca566_u0<=1'h0;
else reg_7d7ca566_u0<=reg_2901482a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_737da366_u0<=1'h0;
else reg_737da366_u0<=reg_039aa343_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5e49b654_u0<=1'h0;
else reg_5e49b654_u0<=reg_60f8cda6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1b5b6b45_u0<=1'h0;
else reg_1b5b6b45_u0<=reg_2a6d54d5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_619c0582_u0<=1'h0;
else reg_619c0582_u0<=reg_062cdef7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1bf28bed_u0<=1'h0;
else reg_1bf28bed_u0<=reg_586b6c26_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1b5b6b45_result_delayed_u0<=1'h0;
else reg_1b5b6b45_result_delayed_u0<=reg_1b5b6b45_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1dc331e7_u0<=1'h0;
else reg_1dc331e7_u0<=reg_42c05205_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_718f51a9_u0<=1'h0;
else reg_718f51a9_u0<=reg_11cd6f36_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1b10bf37_u0<=1'h0;
else reg_1b10bf37_u0<=reg_0924240b_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_44949cbe_u0<=1'h0;
else reg_44949cbe_u0<=reg_09f461a1_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3c729058_u0<=1'h0;
else reg_3c729058_u0<=reg_3736a309_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_69b415a1_result_delayed_u0<=1'h0;
else reg_69b415a1_result_delayed_u0<=reg_69b415a1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_41edcddd_u0<=1'h0;
else reg_41edcddd_u0<=reg_3126cd62_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4ef81ecb_u0<=1'h0;
else reg_4ef81ecb_u0<=reg_2499b3e8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_55610952_u0<=1'h0;
else reg_55610952_u0<=reg_737be907_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_29f9ddea_result_delayed_u0<=1'h0;
else reg_29f9ddea_result_delayed_u0<=reg_29f9ddea_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_787cb445_u0<=1'h0;
else reg_787cb445_u0<=reg_6a945bc0_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5d8aa5b1_u0<=1'h0;
else reg_5d8aa5b1_u0<=reg_2dc36fb8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_632eeb10_u0<=1'h0;
else reg_632eeb10_u0<=reg_7d7ca566_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3736a309_u0<=1'h0;
else reg_3736a309_u0<=reg_4b05af4d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_62a002e4_u0<=1'h0;
else reg_62a002e4_u0<=reg_2ce4bd89_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3126cd62_u0<=1'h0;
else reg_3126cd62_u0<=reg_4a825e39_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5d242960_u0<=1'h0;
else reg_5d242960_u0<=reg_33a8b808_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4b05af4d_u0<=1'h0;
else reg_4b05af4d_u0<=reg_5d8aa5b1_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_586b6c26_u0<=1'h0;
else reg_586b6c26_u0<=reg_51004f81_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3fddb792_u0<=1'h0;
else reg_3fddb792_u0<=reg_0993b092_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_41edcddd_result_delayed_u0<=1'h0;
else reg_41edcddd_result_delayed_u0<=reg_41edcddd_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2ddf258d_u0<=1'h0;
else reg_2ddf258d_u0<=reg_28e17c75_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1af85aaa_u0<=1'h0;
else reg_1af85aaa_u0<=reg_46946686_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_09f461a1_u0<=1'h0;
else reg_09f461a1_u0<=reg_190e5b6d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_25cb699d_u0<=1'h0;
else reg_25cb699d_u0<=reg_1b10bf37_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1f76a321_u0<=1'h0;
else reg_1f76a321_u0<=reg_62a002e4_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6768af3f_u0<=1'h0;
else reg_6768af3f_u0<=reg_67de13aa_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2c47481f_u0<=1'h0;
else reg_2c47481f_u0<=reg_4a991a10_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_04a958f3_u0<=1'h0;
else reg_04a958f3_u0<=reg_63cbe06a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7b1fd745_u0<=1'h0;
else reg_7b1fd745_u0<=reg_1dbaf9d0_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0ac26e9c_u0<=1'h0;
else reg_0ac26e9c_u0<=reg_633a5b40_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1febb7b4_u0<=1'h0;
else reg_1febb7b4_u0<=reg_392f0d9b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_47f4e3ab_u0<=1'h0;
else reg_47f4e3ab_u0<=reg_77462671_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1ed112b0_u0<=1'h0;
else reg_1ed112b0_u0<=reg_0ac6524e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7624ba47_u0<=1'h0;
else reg_7624ba47_u0<=reg_05b504f5_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_47e56b81_u0<=1'h0;
else reg_47e56b81_u0<=and_delayed_u239;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2c204028_result_delayed_u0<=1'h0;
else reg_2c204028_result_delayed_u0<=reg_2c204028_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3765130d_u0<=1'h0;
else reg_3765130d_u0<=reg_4874c2bd_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_47c77fae_u0<=1'h0;
else reg_47c77fae_u0<=reg_3a62176b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1dbaf9d0_u0<=1'h0;
else reg_1dbaf9d0_u0<=reg_73ced32a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_79ff2594_u0<=1'h0;
else reg_79ff2594_u0<=reg_3912a11e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_549798fc_u0<=1'h0;
else reg_549798fc_u0<=reg_2d083c40_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7834905a_u0<=1'h0;
else reg_7834905a_u0<=reg_7a5ce622_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_408e14fc_u0<=1'h0;
else reg_408e14fc_u0<=reg_32d59a7c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a2b825f_u0<=1'h0;
else reg_7a2b825f_u0<=reg_4c4df618_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_67de13aa_u0<=1'h0;
else reg_67de13aa_u0<=reg_45535925_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_45535925_u0<=1'h0;
else reg_45535925_u0<=reg_2d501b7f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_28e2989b_u0<=1'h0;
else reg_28e2989b_u0<=reg_3afa1e08_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_633a5b40_u0<=1'h0;
else reg_633a5b40_u0<=reg_1742dbd1_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3471a47b_result_delayed_u0<=1'h0;
else reg_3471a47b_result_delayed_u0<=reg_3471a47b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3912a11e_result_delayed_u0<=1'h0;
else reg_3912a11e_result_delayed_u0<=reg_3912a11e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a5ce622_u0<=1'h0;
else reg_7a5ce622_u0<=reg_07488981_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5b32ffb2_u0<=1'h0;
else reg_5b32ffb2_u0<=reg_408e14fc_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_71b3a931_u0<=1'h0;
else reg_71b3a931_u0<=reg_65dbefa4_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_23c90b4d_u0<=1'h0;
else reg_23c90b4d_u0<=reg_3a1feec1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_19b1e534_u0<=1'h0;
else reg_19b1e534_u0<=reg_1b2287cc_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_18b39c34_u0<=1'h0;
else reg_18b39c34_u0<=reg_3d2ae849_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0ac6524e_u0<=1'h0;
else reg_0ac6524e_u0<=reg_5236af83_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4a991a10_u0<=1'h0;
else reg_4a991a10_u0<=reg_3b2ea222_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2bd5f75e_u0<=1'h0;
else reg_2bd5f75e_u0<=reg_5e962850_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_005750dc_u0<=1'h0;
else reg_005750dc_u0<=reg_3471a47b_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_67de13aa_result_delayed_u0<=1'h0;
else reg_67de13aa_result_delayed_u0<=reg_67de13aa_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_029c8613_u0<=1'h0;
else reg_029c8613_u0<=reg_4da6e166_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_039f5f0f_u0<=1'h0;
else reg_039f5f0f_u0<=reg_3052e1e7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_31ec057e_u0<=1'h0;
else reg_31ec057e_u0<=reg_28bd586b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1742dbd1_u0<=1'h0;
else reg_1742dbd1_u0<=reg_4c87c45c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_28e17c75_u0<=1'h0;
else reg_28e17c75_u0<=reg_18b39c34_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7fe56773_u0<=1'h0;
else reg_7fe56773_u0<=reg_12299b2b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7dcd9154_u0<=1'h0;
else reg_7dcd9154_u0<=reg_55610952_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_15d1894b_u0<=1'h0;
else reg_15d1894b_u0<=reg_719347fd_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_66fd0261_u0<=1'h0;
else reg_66fd0261_u0<=reg_3de6494b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_25cb699d_result_delayed_u0<=1'h0;
else reg_25cb699d_result_delayed_u0<=reg_25cb699d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_408e14fc_result_delayed_u0<=1'h0;
else reg_408e14fc_result_delayed_u0<=reg_408e14fc_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1dbaf9d0_result_delayed_u0<=1'h0;
else reg_1dbaf9d0_result_delayed_u0<=reg_1dbaf9d0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_34478ce7_u0<=1'h0;
else reg_34478ce7_u0<=reg_1ed112b0_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7b86d327_u0<=1'h0;
else reg_7b86d327_u0<=reg_1b5b6b45_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_44949cbe_result_delayed_u0<=1'h0;
else reg_44949cbe_result_delayed_u0<=reg_44949cbe_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_446bb0cd_u0<=1'h0;
else reg_446bb0cd_u0<=reg_3d4fe5be_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_449ea438_u0<=1'h0;
else reg_449ea438_u0<=reg_1a8ce0d2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_32d59a7c_u0<=1'h0;
else reg_32d59a7c_u0<=reg_50e10aad_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5fce0764_u0<=1'h0;
else reg_5fce0764_u0<=reg_1b78238d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7432b099_u0<=1'h0;
else reg_7432b099_u0<=reg_1cb40934_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3471a47b_result_delayed_result_delayed_u0<=1'h0;
else reg_3471a47b_result_delayed_result_delayed_u0<=reg_3471a47b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3de6494b_u0<=1'h0;
else reg_3de6494b_u0<=reg_2e453868_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_527dd6cc_u0<=1'h0;
else reg_527dd6cc_u0<=reg_3765130d_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6fd8576b_u0<=1'h0;
else reg_6fd8576b_u0<=reg_446bb0cd_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_392f0d9b_u0<=1'h0;
else reg_392f0d9b_u0<=reg_44949cbe_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4a825e39_u0<=1'h0;
else reg_4a825e39_u0<=reg_527dd6cc_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2c204028_result_delayed_result_delayed_u0<=1'h0;
else reg_2c204028_result_delayed_result_delayed_u0<=reg_2c204028_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4da6e166_u0<=1'h0;
else reg_4da6e166_u0<=reg_69b415a1_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_713e21fb_u0<=1'h0;
else reg_713e21fb_u0<=reg_44b53de6_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5d8aa5b1_result_delayed_u0<=1'h0;
else reg_5d8aa5b1_result_delayed_u0<=reg_5d8aa5b1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_42c05205_u0<=1'h0;
else reg_42c05205_u0<=reg_7fca9f36_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_449ea438_result_delayed_u0<=1'h0;
else reg_449ea438_result_delayed_u0<=reg_449ea438_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_11f3093e_u0<=1'h0;
else reg_11f3093e_u0<=reg_1f76a321_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4c2ecce3_u0<=1'h0;
else reg_4c2ecce3_u0<=and_u3612_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_350541ca_u0<=1'h0;
else reg_350541ca_u0<=reg_08ab9607_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7cb11462_u0<=1'h0;
else reg_7cb11462_u0<=reg_568a337f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_45a71573_u0<=1'h0;
else reg_45a71573_u0<=reg_7fa5f2e1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_28bd586b_u0<=1'h0;
else reg_28bd586b_u0<=reg_1f3d20af_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_44949cbe_result_delayed_result_delayed_u0<=1'h0;
else reg_44949cbe_result_delayed_result_delayed_u0<=reg_44949cbe_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_368fce58_u0<=1'h0;
else reg_368fce58_u0<=reg_5cd550db_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_039aa343_u0<=1'h0;
else reg_039aa343_u0<=reg_42fabc9d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4c87c45c_u0<=1'h0;
else reg_4c87c45c_u0<=reg_71134e38_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_062cdef7_u0<=1'h0;
else reg_062cdef7_u0<=reg_713e21fb_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3a1feec1_u0<=1'h0;
else reg_3a1feec1_u0<=reg_26a95b50_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6f802f62_u0<=1'h0;
else reg_6f802f62_u0<=reg_15d1894b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_73ced32a_u0<=1'h0;
else reg_73ced32a_u0<=reg_0f03e5b9_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1cc24c27_u0<=1'h0;
else reg_1cc24c27_u0<=reg_1611b424_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7b9f9b79_u0<=1'h0;
else reg_7b9f9b79_u0<=reg_632eeb10_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2ae45e03_u0<=1'h0;
else reg_2ae45e03_u0<=reg_3fddb792_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1b2287cc_u0<=1'h0;
else reg_1b2287cc_u0<=reg_41edcddd_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3d4fe5be_u0<=1'h0;
else reg_3d4fe5be_u0<=reg_04a958f3_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3afa1e08_u0<=1'h0;
else reg_3afa1e08_u0<=reg_602c59ab_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1ba0d353_u0<=1'h0;
else reg_1ba0d353_u0<=reg_0525586a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1b78238d_u0<=1'h0;
else reg_1b78238d_u0<=reg_49656763_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2632face_u0<=1'h0;
else reg_2632face_u0<=reg_1bf28bed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7fca9f36_u0<=1'h0;
else reg_7fca9f36_u0<=reg_0b45c90a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7dd95126_u0<=1'h0;
else reg_7dd95126_u0<=reg_4ff65e34_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0993b092_u0<=1'h0;
else reg_0993b092_u0<=reg_6e167f08_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_12299b2b_u0<=1'h0;
else reg_12299b2b_u0<=reg_1324a63d_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7ce161e2_u0<=1'h0;
else reg_7ce161e2_u0<=reg_71d3e4cd_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7ce161e2_result_delayed_u0<=1'h0;
else reg_7ce161e2_result_delayed_u0<=reg_7ce161e2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3a62176b_u0<=1'h0;
else reg_3a62176b_u0<=reg_30e129c3_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_029c8613_result_delayed_u0<=1'h0;
else reg_029c8613_result_delayed_u0<=reg_029c8613_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01539059_u0<=1'h0;
else reg_01539059_u0<=reg_13ea2607_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4bc316c8_u0<=1'h0;
else reg_4bc316c8_u0<=reg_6f802f62_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0af8dff3_u0<=1'h0;
else reg_0af8dff3_u0<=reg_61ecb46b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_69ccc0c7_u0<=1'h0;
else reg_69ccc0c7_u0<=reg_3c844144_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7432b099_result_delayed_u0<=1'h0;
else reg_7432b099_result_delayed_u0<=reg_7432b099_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3b2ea222_u0<=1'h0;
else reg_3b2ea222_u0<=reg_69f58839_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5792329f_u0<=1'h0;
else reg_5792329f_u0<=reg_7b86d327_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_46946686_result_delayed_u0<=1'h0;
else reg_46946686_result_delayed_u0<=reg_46946686_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_67e61ef6_u0<=1'h0;
else reg_67e61ef6_u0<=reg_2fe53643_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3471a47b_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_3471a47b_result_delayed_result_delayed_result_delayed_u0<=reg_3471a47b_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1b5b6b45_result_delayed_result_delayed_u0<=1'h0;
else reg_1b5b6b45_result_delayed_result_delayed_u0<=reg_1b5b6b45_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_70705567_u0<=1'h0;
else reg_70705567_u0<=reg_0188e8a7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1324a63d_u0<=1'h0;
else reg_1324a63d_u0<=reg_0ac26e9c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2ae45e03_result_delayed_u0<=1'h0;
else reg_2ae45e03_result_delayed_u0<=reg_2ae45e03_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3afa1e08_result_delayed_u0<=1'h0;
else reg_3afa1e08_result_delayed_u0<=reg_3afa1e08_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_71d3e4cd_u0<=1'h0;
else reg_71d3e4cd_u0<=reg_3db3d453_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6e167f08_u0<=1'h0;
else reg_6e167f08_u0<=reg_6a83a8be_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4012210d_u0<=1'h0;
else reg_4012210d_u0<=reg_7a349f51_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0127d038_u0<=1'h0;
else reg_0127d038_u0<=reg_43dd6207_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_30e129c3_u0<=1'h0;
else reg_30e129c3_u0<=reg_7624ba47_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2b525e7b_u0<=1'h0;
else reg_2b525e7b_u0<=reg_351e991f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_134a2263_u0<=1'h0;
else reg_134a2263_u0<=reg_74967c94_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_70705567_result_delayed_u0<=1'h0;
else reg_70705567_result_delayed_u0<=reg_70705567_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2901482a_u0<=1'h0;
else reg_2901482a_u0<=reg_1554b782_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0924240b_u0<=1'h0;
else reg_0924240b_u0<=reg_2632face_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0188e8a7_u0<=1'h0;
else reg_0188e8a7_u0<=reg_3c729058_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3afa1e08_result_delayed_result_delayed_u0<=1'h0;
else reg_3afa1e08_result_delayed_result_delayed_u0<=reg_3afa1e08_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_63aaa29e_u0<=1'h0;
else reg_63aaa29e_u0<=reg_0f0fdd38_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_77462671_u0<=1'h0;
else reg_77462671_u0<=reg_5d242960_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_408e14fc_result_delayed_result_delayed_u0<=1'h0;
else reg_408e14fc_result_delayed_result_delayed_u0<=reg_408e14fc_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_446bb0cd_result_delayed_u0<=1'h0;
else reg_446bb0cd_result_delayed_u0<=reg_446bb0cd_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_527dd6cc_result_delayed_u0<=1'h0;
else reg_527dd6cc_result_delayed_u0<=reg_527dd6cc_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_05b504f5_u0<=1'h0;
else reg_05b504f5_u0<=reg_2377f2f2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7b991f92_result_delayed_u0<=1'h0;
else reg_7b991f92_result_delayed_u0<=reg_7b991f92_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7fa5f2e1_u0<=1'h0;
else reg_7fa5f2e1_u0<=reg_622e780a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5fc7b281_u0<=1'h0;
else reg_5fc7b281_u0<=reg_1af85aaa_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_08cf2d88_u0<=1'h0;
else reg_08cf2d88_u0<=reg_4ef81ecb_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2d083c40_u0<=1'h0;
else reg_2d083c40_u0<=reg_350541ca_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_62aecfe4_u0<=1'h0;
else reg_62aecfe4_u0<=reg_010e94b1_result_delayed_u0;
end
assign and_u3611_u0=and_u3606_u0&and_u3613_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_449ea438_result_delayed_result_delayed_u0<=1'h0;
else reg_449ea438_result_delayed_result_delayed_u0<=reg_449ea438_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0525586a_u0<=1'h0;
else reg_0525586a_u0<=reg_28e2989b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_25cb699d_result_delayed_result_delayed_u0<=1'h0;
else reg_25cb699d_result_delayed_result_delayed_u0<=reg_25cb699d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4f8742d5_u0<=1'h0;
else reg_4f8742d5_u0<=reg_6a850ff6_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_350541ca_result_delayed_u0<=1'h0;
else reg_350541ca_result_delayed_u0<=reg_350541ca_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_44b53de6_u0<=1'h0;
else reg_44b53de6_u0<=reg_2b525e7b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6a945bc0_u0<=1'h0;
else reg_6a945bc0_u0<=reg_29f9ddea_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5d8aa5b1_result_delayed_result_delayed_u0<=1'h0;
else reg_5d8aa5b1_result_delayed_result_delayed_u0<=reg_5d8aa5b1_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4b05af4d_result_delayed_u0<=1'h0;
else reg_4b05af4d_result_delayed_u0<=reg_4b05af4d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_619c0582_result_delayed_u0<=1'h0;
else reg_619c0582_result_delayed_u0<=reg_619c0582_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_60f8cda6_u0<=1'h0;
else reg_60f8cda6_u0<=reg_7ee659a2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1801415e_u0<=1'h0;
else reg_1801415e_u0<=reg_5b32ffb2_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1ec2c3a2_u0<=1'h0;
else reg_1ec2c3a2_u0<=reg_5e49b654_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_74967c94_result_delayed_result_delayed_u0<=1'h0;
else reg_74967c94_result_delayed_result_delayed_u0<=reg_74967c94_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_12bc27dd_u0<=1'h0;
else reg_12bc27dd_u0<=reg_70705567_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3d2ae849_u0<=1'h0;
else reg_3d2ae849_u0<=reg_57b957bf_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a349f51_u0<=1'h0;
else reg_7a349f51_u0<=reg_697bf970_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_62aecfe4_result_delayed_u0<=1'h0;
else reg_62aecfe4_result_delayed_u0<=reg_62aecfe4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_47e56b81_result_delayed_u0<=1'h0;
else reg_47e56b81_result_delayed_u0<=reg_47e56b81_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0ac26e9c_result_delayed_u0<=1'h0;
else reg_0ac26e9c_result_delayed_u0<=reg_0ac26e9c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2ce4bd89_u0<=1'h0;
else reg_2ce4bd89_u0<=reg_549798fc_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_27d7caa5_u0<=1'h0;
else reg_27d7caa5_u0<=reg_1dca001c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6a850ff6_u0<=1'h0;
else reg_6a850ff6_u0<=reg_51cd934d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_12bc27dd_result_delayed_u0<=1'h0;
else reg_12bc27dd_result_delayed_u0<=reg_12bc27dd_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7f9742e2_u0<=1'h0;
else reg_7f9742e2_u0<=reg_3b9cf399_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_719ae8ef_u0<=1'h0;
else reg_719ae8ef_u0<=reg_193758c8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6efe4388_u0<=1'h0;
else reg_6efe4388_u0<=reg_0af8dff3_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1801415e_result_delayed_u0<=1'h0;
else reg_1801415e_result_delayed_u0<=reg_1801415e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1cb40934_u0<=1'h0;
else reg_1cb40934_u0<=reg_582b1a27_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_351e991f_result_delayed_u0<=1'h0;
else reg_351e991f_result_delayed_u0<=reg_351e991f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_10d31157_u0<=1'h0;
else reg_10d31157_u0<=reg_7fe56773_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2377f2f2_u0<=1'h0;
else reg_2377f2f2_u0<=reg_47e56b81_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_61ecb46b_u0<=1'h0;
else reg_61ecb46b_u0<=reg_3ef9b436_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_602c59ab_u0<=1'h0;
else reg_602c59ab_u0<=reg_049d62ec_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_41edcddd_result_delayed_result_delayed_u0<=1'h0;
else reg_41edcddd_result_delayed_result_delayed_u0<=reg_41edcddd_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_54ab7523_u0<=1'h0;
else reg_54ab7523_u0<=reg_23c90b4d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_385515de_u0<=1'h0;
else reg_385515de_u0<=reg_7b991f92_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6a945bc0_result_delayed_u0<=1'h0;
else reg_6a945bc0_result_delayed_u0<=reg_6a945bc0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_03b7ae24_u0<=1'h0;
else reg_03b7ae24_u0<=reg_1ba0d353_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3765130d_result_delayed_u0<=1'h0;
else reg_3765130d_result_delayed_u0<=reg_3765130d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2b525e7b_result_delayed_u0<=1'h0;
else reg_2b525e7b_result_delayed_u0<=reg_2b525e7b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7121f4b8_u0<=1'h0;
else reg_7121f4b8_u0<=reg_4650dc26_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_52798be3_u0<=1'h0;
else reg_52798be3_u0<=reg_1130ef58_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5e49b654_result_delayed_u0<=1'h0;
else reg_5e49b654_result_delayed_u0<=reg_5e49b654_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2fe53643_u0<=1'h0;
else reg_2fe53643_u0<=reg_633a799d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2c47481f_result_delayed_u0<=1'h0;
else reg_2c47481f_result_delayed_u0<=reg_2c47481f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_37b15a18_u0<=1'h0;
else reg_37b15a18_u0<=reg_60d46663_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6efe4388_result_delayed_u0<=1'h0;
else reg_6efe4388_result_delayed_u0<=reg_6efe4388_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3052e1e7_u0<=1'h0;
else reg_3052e1e7_u0<=reg_52798be3_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5236af83_u0<=1'h0;
else reg_5236af83_u0<=reg_039f5f0f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7b1fd745_result_delayed_u0<=1'h0;
else reg_7b1fd745_result_delayed_u0<=reg_7b1fd745_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_010e94b1_u0<=1'h0;
else reg_010e94b1_u0<=reg_7b1fd745_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3c844144_u0<=1'h0;
else reg_3c844144_u0<=reg_2ded6345_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0af8dff3_result_delayed_u0<=1'h0;
else reg_0af8dff3_result_delayed_u0<=reg_0af8dff3_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4ff65e34_u0<=1'h0;
else reg_4ff65e34_u0<=reg_1dc331e7_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_69b415a1_result_delayed_result_delayed_u0<=1'h0;
else reg_69b415a1_result_delayed_result_delayed_u0<=reg_69b415a1_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_69f58839_u0<=1'h0;
else reg_69f58839_u0<=reg_47f4e3ab_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_719ae8ef_result_delayed_u0<=1'h0;
else reg_719ae8ef_result_delayed_u0<=reg_719ae8ef_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1ed112b0_result_delayed_u0<=1'h0;
else reg_1ed112b0_result_delayed_u0<=reg_1ed112b0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_16e37f2c_u0<=1'h0;
else reg_16e37f2c_u0<=reg_1cc24c27_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3fddb792_result_delayed_u0<=1'h0;
else reg_3fddb792_result_delayed_u0<=reg_3fddb792_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1dca001c_u0<=1'h0;
else reg_1dca001c_u0<=reg_15fe439b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_08cf2d88_result_delayed_u0<=1'h0;
else reg_08cf2d88_result_delayed_u0<=reg_08cf2d88_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_43dd6207_u0<=1'h0;
else reg_43dd6207_u0<=reg_4012210d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0bd5de0a_u0<=1'h0;
else reg_0bd5de0a_u0<=reg_092d4389_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3db3d453_u0<=1'h0;
else reg_3db3d453_u0<=reg_17bf09db_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3765130d_result_delayed_result_delayed_u0<=1'h0;
else reg_3765130d_result_delayed_result_delayed_u0<=reg_3765130d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_713e21fb_result_delayed_u0<=1'h0;
else reg_713e21fb_result_delayed_u0<=reg_713e21fb_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1dbaf9d0_result_delayed_result_delayed_u0<=1'h0;
else reg_1dbaf9d0_result_delayed_result_delayed_u0<=reg_1dbaf9d0_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_13ea2607_u0<=1'h0;
else reg_13ea2607_u0<=reg_7dd95126_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0924240b_result_delayed_u0<=1'h0;
else reg_0924240b_result_delayed_u0<=reg_0924240b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3c729058_result_delayed_u0<=1'h0;
else reg_3c729058_result_delayed_u0<=reg_3c729058_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u239<=1'h0;
else and_delayed_u239<=and_u3611_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_005750dc_result_delayed_u0<=1'h0;
else reg_005750dc_result_delayed_u0<=reg_005750dc_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_568a337f_u0<=1'h0;
else reg_568a337f_u0<=reg_3c1b12e8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1742dbd1_result_delayed_u0<=1'h0;
else reg_1742dbd1_result_delayed_u0<=reg_1742dbd1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_26a95b50_u0<=1'h0;
else reg_26a95b50_u0<=reg_1801415e_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2fbb9e45_u0<=1'h0;
else reg_2fbb9e45_u0<=reg_69ccc0c7_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_193758c8_u0<=1'h0;
else reg_193758c8_u0<=reg_40f3fed8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_713c4f38_u0<=1'h0;
else reg_713c4f38_u0<=reg_787cb445_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_49656763_u0<=1'h0;
else reg_49656763_u0<=reg_2c47481f_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6bfaddf3_u0<=1'h0;
else reg_6bfaddf3_u0<=reg_25cb699d_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1cc24c27_result_delayed_u0<=1'h0;
else reg_1cc24c27_result_delayed_u0<=reg_1cc24c27_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_582b1a27_u0<=1'h0;
else reg_582b1a27_u0<=reg_385515de_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_527dd6cc_result_delayed_result_delayed_u0<=1'h0;
else reg_527dd6cc_result_delayed_result_delayed_u0<=reg_527dd6cc_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_787cb445_result_delayed_u0<=1'h0;
else reg_787cb445_result_delayed_u0<=reg_787cb445_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01539059_result_delayed_u0<=1'h0;
else reg_01539059_result_delayed_u0<=reg_01539059_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_622e780a_u0<=1'h0;
else reg_622e780a_u0<=reg_6efe4388_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5cd550db_result_delayed_u0<=1'h0;
else reg_5cd550db_result_delayed_u0<=reg_5cd550db_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_40f3fed8_u0<=1'h0;
else reg_40f3fed8_u0<=reg_449ea438_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2e453868_u0<=1'h0;
else reg_2e453868_u0<=reg_62aecfe4_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2d501b7f_u0<=1'h0;
else reg_2d501b7f_u0<=reg_63aaa29e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_449ea438_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_449ea438_result_delayed_result_delayed_result_delayed_u0<=reg_449ea438_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1611b424_u0<=1'h0;
else reg_1611b424_u0<=reg_1ec2c3a2_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0f0fdd38_u0<=1'h0;
else reg_0f0fdd38_u0<=reg_16e37f2c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_582b1a27_result_delayed_u0<=1'h0;
else reg_582b1a27_result_delayed_u0<=reg_582b1a27_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1b10bf37_result_delayed_u0<=1'h0;
else reg_1b10bf37_result_delayed_u0<=reg_1b10bf37_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6a83a8be_u0<=1'h0;
else reg_6a83a8be_u0<=reg_617de3bd_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_713e21fb_result_delayed_result_delayed_u0<=1'h0;
else reg_713e21fb_result_delayed_result_delayed_u0<=reg_713e21fb_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_37b15a18_result_delayed_u0<=1'h0;
else reg_37b15a18_result_delayed_u0<=reg_37b15a18_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_12e4f0a0_u0<=1'h0;
else reg_12e4f0a0_u0<=reg_286c1a08_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_29f9ddea_result_delayed_result_delayed_u0<=1'h0;
else reg_29f9ddea_result_delayed_result_delayed_u0<=reg_29f9ddea_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_787cb445_result_delayed_result_delayed_u0<=1'h0;
else reg_787cb445_result_delayed_result_delayed_u0<=reg_787cb445_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_50e10aad_u0<=1'h0;
else reg_50e10aad_u0<=reg_005750dc_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0b45c90a_u0<=1'h0;
else reg_0b45c90a_u0<=reg_0224b0d4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0820ce74_u0<=1'h0;
else reg_0820ce74_u0<=reg_5dc782c5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4c4df618_u0<=1'h0;
else reg_4c4df618_u0<=reg_5792329f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_55610952_result_delayed_u0<=1'h0;
else reg_55610952_result_delayed_u0<=reg_55610952_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7b1fd745_result_delayed_result_delayed_u0<=1'h0;
else reg_7b1fd745_result_delayed_result_delayed_u0<=reg_7b1fd745_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_79ff2594_result_delayed_u0<=1'h0;
else reg_79ff2594_result_delayed_u0<=reg_79ff2594_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1a8ce0d2_u0<=1'h0;
else reg_1a8ce0d2_u0<=reg_713c4f38_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_190e5b6d_u0<=1'h0;
else reg_190e5b6d_u0<=reg_45a71573_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_286c1a08_u0<=1'h0;
else reg_286c1a08_u0<=reg_0820ce74_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_17bf09db_u0<=1'h0;
else reg_17bf09db_u0<=reg_27d7caa5_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_15fe439b_u0<=1'h0;
else reg_15fe439b_u0<=reg_36c619e0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7624ba47_result_delayed_u0<=1'h0;
else reg_7624ba47_result_delayed_u0<=reg_7624ba47_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_42fabc9d_u0<=1'h0;
else reg_42fabc9d_u0<=reg_4bc316c8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1130ef58_u0<=1'h0;
else reg_1130ef58_u0<=reg_7ce161e2_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6a83a8be_result_delayed_u0<=1'h0;
else reg_6a83a8be_result_delayed_u0<=reg_6a83a8be_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_47f4e3ab_result_delayed_u0<=1'h0;
else reg_47f4e3ab_result_delayed_u0<=reg_47f4e3ab_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_719347fd_u0<=1'h0;
else reg_719347fd_u0<=reg_6a948183_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6a945bc0_result_delayed_result_delayed_u0<=1'h0;
else reg_6a945bc0_result_delayed_result_delayed_u0<=reg_6a945bc0_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a2b825f_result_delayed_u0<=1'h0;
else reg_7a2b825f_result_delayed_u0<=reg_7a2b825f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_049d62ec_u0<=1'h0;
else reg_049d62ec_u0<=reg_66fd0261_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1795d1e7_u0<=1'h0;
else reg_1795d1e7_u0<=reg_486de694_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_62a002e4_result_delayed_u0<=1'h0;
else reg_62a002e4_result_delayed_u0<=reg_62a002e4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4650dc26_u0<=1'h0;
else reg_4650dc26_u0<=reg_67e61ef6_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5b32ffb2_result_delayed_u0<=1'h0;
else reg_5b32ffb2_result_delayed_u0<=reg_5b32ffb2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1f76a321_result_delayed_u0<=1'h0;
else reg_1f76a321_result_delayed_u0<=reg_1f76a321_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2dc36fb8_u0<=1'h0;
else reg_2dc36fb8_u0<=reg_029c8613_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_737be907_u0<=1'h0;
else reg_737be907_u0<=reg_2ae45e03_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_09f461a1_result_delayed_u0<=1'h0;
else reg_09f461a1_result_delayed_u0<=reg_09f461a1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_65dbefa4_u0<=1'h0;
else reg_65dbefa4_u0<=reg_69e5773a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_51cd934d_u0<=1'h0;
else reg_51cd934d_u0<=reg_718f51a9_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_51004f81_u0<=1'h0;
else reg_51004f81_u0<=reg_37d2817c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_69ccc0c7_result_delayed_u0<=1'h0;
else reg_69ccc0c7_result_delayed_u0<=reg_69ccc0c7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0924240b_result_delayed_result_delayed_u0<=1'h0;
else reg_0924240b_result_delayed_result_delayed_u0<=reg_0924240b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_549798fc_result_delayed_u0<=1'h0;
else reg_549798fc_result_delayed_u0<=reg_549798fc_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_67e61ef6_result_delayed_u0<=1'h0;
else reg_67e61ef6_result_delayed_u0<=reg_67e61ef6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_69f58839_result_delayed_u0<=1'h0;
else reg_69f58839_result_delayed_u0<=reg_69f58839_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3d2ae849_result_delayed_u0<=1'h0;
else reg_3d2ae849_result_delayed_u0<=reg_3d2ae849_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1b5b6b45_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_1b5b6b45_result_delayed_result_delayed_result_delayed_u0<=reg_1b5b6b45_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_41edcddd_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_41edcddd_result_delayed_result_delayed_result_delayed_u0<=reg_41edcddd_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1dbaf9d0_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_1dbaf9d0_result_delayed_result_delayed_result_delayed_u0<=reg_1dbaf9d0_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6fd8576b_result_delayed_u0<=1'h0;
else reg_6fd8576b_result_delayed_u0<=reg_6fd8576b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_190e5b6d_result_delayed_u0<=1'h0;
else reg_190e5b6d_result_delayed_u0<=reg_190e5b6d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_26a95b50_result_delayed_u0<=1'h0;
else reg_26a95b50_result_delayed_u0<=reg_26a95b50_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_57b957bf_result_delayed_u0<=1'h0;
else reg_57b957bf_result_delayed_u0<=reg_57b957bf_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_549798fc_result_delayed_result_delayed_u0<=1'h0;
else reg_549798fc_result_delayed_result_delayed_u0<=reg_549798fc_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_44b53de6_result_delayed_u0<=1'h0;
else reg_44b53de6_result_delayed_u0<=reg_44b53de6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2fe53643_result_delayed_u0<=1'h0;
else reg_2fe53643_result_delayed_u0<=reg_2fe53643_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_010e94b1_result_delayed_u0<=1'h0;
else reg_010e94b1_result_delayed_u0<=reg_010e94b1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7ce161e2_result_delayed_result_delayed_u0<=1'h0;
else reg_7ce161e2_result_delayed_result_delayed_u0<=reg_7ce161e2_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_092d4389_u0<=1'h0;
else reg_092d4389_u0<=reg_57e6dcb6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7cb11462_result_delayed_u0<=1'h0;
else reg_7cb11462_result_delayed_u0<=reg_7cb11462_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_633a799d_u0<=1'h0;
else reg_633a799d_u0<=reg_7f9742e2_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2ded6345_u0<=1'h0;
else reg_2ded6345_u0<=reg_5fc7b281_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0db7cb1d_u0<=1'h0;
else reg_0db7cb1d_u0<=reg_54ab7523_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7fe56773_result_delayed_u0<=1'h0;
else reg_7fe56773_result_delayed_u0<=reg_7fe56773_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_08ab9607_u0<=1'h0;
else reg_08ab9607_u0<=reg_2ddf258d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_37d2817c_u0<=1'h0;
else reg_37d2817c_u0<=reg_47c77fae_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_12247897_u0<=1'h0;
else reg_12247897_u0<=reg_719ae8ef_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4c4df618_result_delayed_u0<=1'h0;
else reg_4c4df618_result_delayed_u0<=reg_4c4df618_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_67e61ef6_result_delayed_result_delayed_u0<=1'h0;
else reg_67e61ef6_result_delayed_result_delayed_u0<=reg_67e61ef6_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_60d46663_u0<=1'h0;
else reg_60d46663_u0<=reg_072dadc1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2a6d54d5_u0<=1'h0;
else reg_2a6d54d5_u0<=reg_79ff2594_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0f03e5b9_u0<=1'h0;
else reg_0f03e5b9_u0<=reg_12247897_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5792329f_result_delayed_u0<=1'h0;
else reg_5792329f_result_delayed_u0<=reg_5792329f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2632face_result_delayed_u0<=1'h0;
else reg_2632face_result_delayed_u0<=reg_2632face_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2bd5f75e_result_delayed_u0<=1'h0;
else reg_2bd5f75e_result_delayed_u0<=reg_2bd5f75e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_617de3bd_u0<=1'h0;
else reg_617de3bd_u0<=reg_2fbb9e45_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_26a95b50_result_delayed_result_delayed_u0<=1'h0;
else reg_26a95b50_result_delayed_result_delayed_u0<=reg_26a95b50_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6f802f62_result_delayed_u0<=1'h0;
else reg_6f802f62_result_delayed_u0<=reg_6f802f62_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_15fe439b_result_delayed_u0<=1'h0;
else reg_15fe439b_result_delayed_u0<=reg_15fe439b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0ac6524e_result_delayed_u0<=1'h0;
else reg_0ac6524e_result_delayed_u0<=reg_0ac6524e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5e962850_u0<=1'h0;
else reg_5e962850_u0<=reg_31ec057e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4012210d_result_delayed_u0<=1'h0;
else reg_4012210d_result_delayed_u0<=reg_4012210d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_07488981_u0<=1'h0;
else reg_07488981_u0<=reg_7121f4b8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4874c2bd_u0<=1'h0;
else reg_4874c2bd_u0<=reg_08cf2d88_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_582b1a27_result_delayed_result_delayed_u0<=1'h0;
else reg_582b1a27_result_delayed_result_delayed_u0<=reg_582b1a27_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0127d038_result_delayed_u0<=1'h0;
else reg_0127d038_result_delayed_u0<=reg_0127d038_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3ef9b436_u0<=1'h0;
else reg_3ef9b436_u0<=reg_34478ce7_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4f8742d5_result_delayed_u0<=1'h0;
else reg_4f8742d5_result_delayed_u0<=reg_4f8742d5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7121f4b8_result_delayed_u0<=1'h0;
else reg_7121f4b8_result_delayed_u0<=reg_7121f4b8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_27d7caa5_result_delayed_u0<=1'h0;
else reg_27d7caa5_result_delayed_u0<=reg_27d7caa5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_18b39c34_result_delayed_u0<=1'h0;
else reg_18b39c34_result_delayed_u0<=reg_18b39c34_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1554b782_u0<=1'h0;
else reg_1554b782_u0<=reg_46b7b9ba_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2c47481f_result_delayed_result_delayed_u0<=1'h0;
else reg_2c47481f_result_delayed_result_delayed_u0<=reg_2c47481f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1af85aaa_result_delayed_u0<=1'h0;
else reg_1af85aaa_result_delayed_u0<=reg_1af85aaa_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_446bb0cd_result_delayed_result_delayed_u0<=1'h0;
else reg_446bb0cd_result_delayed_result_delayed_u0<=reg_446bb0cd_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_54ab7523_result_delayed_u0<=1'h0;
else reg_54ab7523_result_delayed_u0<=reg_54ab7523_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_69e5773a_u0<=1'h0;
else reg_69e5773a_u0<=reg_7cb11462_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_31ec057e_result_delayed_u0<=1'h0;
else reg_31ec057e_result_delayed_u0<=reg_31ec057e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3471a47b_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_3471a47b_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_3471a47b_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_713e21fb_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_713e21fb_result_delayed_result_delayed_result_delayed_u0<=reg_713e21fb_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_072dadc1_u0<=1'h0;
else reg_072dadc1_u0<=reg_7a2b825f_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_17bf09db_result_delayed_u0<=1'h0;
else reg_17bf09db_result_delayed_u0<=reg_17bf09db_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_70705567_result_delayed_result_delayed_u0<=1'h0;
else reg_70705567_result_delayed_result_delayed_u0<=reg_70705567_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_23c90b4d_result_delayed_u0<=1'h0;
else reg_23c90b4d_result_delayed_u0<=reg_23c90b4d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0224b0d4_u0<=1'h0;
else reg_0224b0d4_u0<=reg_7b9f9b79_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3c1b12e8_u0<=1'h0;
else reg_3c1b12e8_u0<=reg_10d31157_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_27d7caa5_result_delayed_result_delayed_u0<=1'h0;
else reg_27d7caa5_result_delayed_result_delayed_u0<=reg_27d7caa5_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_408e14fc_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_408e14fc_result_delayed_result_delayed_result_delayed_u0<=reg_408e14fc_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_12247897_result_delayed_u0<=1'h0;
else reg_12247897_result_delayed_u0<=reg_12247897_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_486de694_u0<=1'h0;
else reg_486de694_u0<=reg_11f3093e_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_11cd6f36_u0<=1'h0;
else reg_11cd6f36_u0<=reg_37b15a18_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_47f4e3ab_result_delayed_result_delayed_u0<=1'h0;
else reg_47f4e3ab_result_delayed_result_delayed_u0<=reg_47f4e3ab_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_11f3093e_result_delayed_u0<=1'h0;
else reg_11f3093e_result_delayed_u0<=reg_11f3093e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_713c4f38_result_delayed_u0<=1'h0;
else reg_713c4f38_result_delayed_u0<=reg_713c4f38_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5dc782c5_u0<=1'h0;
else reg_5dc782c5_u0<=reg_4f8742d5_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1b2287cc_result_delayed_u0<=1'h0;
else reg_1b2287cc_result_delayed_u0<=reg_1b2287cc_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1dca001c_result_delayed_u0<=1'h0;
else reg_1dca001c_result_delayed_u0<=reg_1dca001c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_46b7b9ba_u0<=1'h0;
else reg_46b7b9ba_u0<=reg_134a2263_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3de6494b_result_delayed_u0<=1'h0;
else reg_3de6494b_result_delayed_u0<=reg_3de6494b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7f9742e2_result_delayed_u0<=1'h0;
else reg_7f9742e2_result_delayed_u0<=reg_7f9742e2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6a948183_u0<=1'h0;
else reg_6a948183_u0<=reg_7834905a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_66fd0261_result_delayed_u0<=1'h0;
else reg_66fd0261_result_delayed_u0<=reg_66fd0261_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5fc7b281_result_delayed_u0<=1'h0;
else reg_5fc7b281_result_delayed_u0<=reg_5fc7b281_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_134a2263_result_delayed_u0<=1'h0;
else reg_134a2263_result_delayed_u0<=reg_134a2263_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a2b825f_result_delayed_result_delayed_u0<=1'h0;
else reg_7a2b825f_result_delayed_result_delayed_u0<=reg_7a2b825f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_36c619e0_u0<=1'h0;
else reg_36c619e0_u0<=reg_51926d82_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_719ae8ef_result_delayed_result_delayed_u0<=1'h0;
else reg_719ae8ef_result_delayed_result_delayed_u0<=reg_719ae8ef_result_delayed_u0;
end
assign and_u3612_u0=and_u3607_u0&and_u3613_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_51926d82_result_delayed_u0<=1'h0;
else reg_51926d82_result_delayed_u0<=reg_51926d82_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_71134e38_u0<=1'h0;
else reg_71134e38_u0<=reg_1febb7b4_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7b86d327_result_delayed_u0<=1'h0;
else reg_7b86d327_result_delayed_u0<=reg_7b86d327_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_28e2989b_result_delayed_u0<=1'h0;
else reg_28e2989b_result_delayed_u0<=reg_28e2989b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_11f3093e_result_delayed_result_delayed_u0<=1'h0;
else reg_11f3093e_result_delayed_result_delayed_u0<=reg_11f3093e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0820ce74_result_delayed_u0<=1'h0;
else reg_0820ce74_result_delayed_u0<=reg_0820ce74_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1554b782_result_delayed_u0<=1'h0;
else reg_1554b782_result_delayed_u0<=reg_1554b782_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_71d3e4cd_result_delayed_u0<=1'h0;
else reg_71d3e4cd_result_delayed_u0<=reg_71d3e4cd_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5d242960_result_delayed_u0<=1'h0;
else reg_5d242960_result_delayed_u0<=reg_5d242960_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_50e10aad_result_delayed_u0<=1'h0;
else reg_50e10aad_result_delayed_u0<=reg_50e10aad_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7ee659a2_u0<=1'h0;
else reg_7ee659a2_u0<=reg_4fad7ce4_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1febb7b4_result_delayed_u0<=1'h0;
else reg_1febb7b4_result_delayed_u0<=reg_1febb7b4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_28e17c75_result_delayed_u0<=1'h0;
else reg_28e17c75_result_delayed_u0<=reg_28e17c75_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4fad7ce4_u0<=1'h0;
else reg_4fad7ce4_u0<=reg_12bc27dd_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_718f51a9_result_delayed_u0<=1'h0;
else reg_718f51a9_result_delayed_u0<=reg_718f51a9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1dc331e7_result_delayed_u0<=1'h0;
else reg_1dc331e7_result_delayed_u0<=reg_1dc331e7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2fbb9e45_result_delayed_u0<=1'h0;
else reg_2fbb9e45_result_delayed_u0<=reg_2fbb9e45_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_47c77fae_result_delayed_u0<=1'h0;
else reg_47c77fae_result_delayed_u0<=reg_47c77fae_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_350541ca_result_delayed_result_delayed_u0<=1'h0;
else reg_350541ca_result_delayed_result_delayed_u0<=reg_350541ca_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1bf28bed_result_delayed_u0<=1'h0;
else reg_1bf28bed_result_delayed_u0<=reg_1bf28bed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_79ff2594_result_delayed_result_delayed_u0<=1'h0;
else reg_79ff2594_result_delayed_result_delayed_u0<=reg_79ff2594_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_57e6dcb6_u0<=1'h0;
else reg_57e6dcb6_u0<=reg_6768af3f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_63aaa29e_result_delayed_u0<=1'h0;
else reg_63aaa29e_result_delayed_u0<=reg_63aaa29e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_05b504f5_result_delayed_u0<=1'h0;
else reg_05b504f5_result_delayed_u0<=reg_05b504f5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2bd5f75e_result_delayed_result_delayed_u0<=1'h0;
else reg_2bd5f75e_result_delayed_result_delayed_u0<=reg_2bd5f75e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_51004f81_result_delayed_u0<=1'h0;
else reg_51004f81_result_delayed_u0<=reg_51004f81_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5d8aa5b1_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_5d8aa5b1_result_delayed_result_delayed_result_delayed_u0<=reg_5d8aa5b1_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_71134e38_result_delayed_u0<=1'h0;
else reg_71134e38_result_delayed_u0<=reg_71134e38_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_385515de_result_delayed_u0<=1'h0;
else reg_385515de_result_delayed_u0<=reg_385515de_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_60d46663_result_delayed_u0<=1'h0;
else reg_60d46663_result_delayed_u0<=reg_60d46663_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_62aecfe4_result_delayed_result_delayed_u0<=1'h0;
else reg_62aecfe4_result_delayed_result_delayed_u0<=reg_62aecfe4_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_08cf2d88_result_delayed_result_delayed_u0<=1'h0;
else reg_08cf2d88_result_delayed_result_delayed_u0<=reg_08cf2d88_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_04a958f3_result_delayed_u0<=1'h0;
else reg_04a958f3_result_delayed_u0<=reg_04a958f3_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_632eeb10_result_delayed_u0<=1'h0;
else reg_632eeb10_result_delayed_u0<=reg_632eeb10_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2ddf258d_result_delayed_u0<=1'h0;
else reg_2ddf258d_result_delayed_u0<=reg_2ddf258d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_549798fc_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_549798fc_result_delayed_result_delayed_result_delayed_u0<=reg_549798fc_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1324a63d_result_delayed_u0<=1'h0;
else reg_1324a63d_result_delayed_u0<=reg_1324a63d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7dd95126_result_delayed_u0<=1'h0;
else reg_7dd95126_result_delayed_u0<=reg_7dd95126_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3a62176b_result_delayed_u0<=1'h0;
else reg_3a62176b_result_delayed_u0<=reg_3a62176b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2499b3e8_u0<=1'h0;
else reg_2499b3e8_u0<=reg_368fce58_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4f8742d5_result_delayed_result_delayed_u0<=1'h0;
else reg_4f8742d5_result_delayed_result_delayed_u0<=reg_4f8742d5_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_15d1894b_result_delayed_u0<=1'h0;
else reg_15d1894b_result_delayed_u0<=reg_15d1894b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_47e56b81_result_delayed_result_delayed_u0<=1'h0;
else reg_47e56b81_result_delayed_result_delayed_u0<=reg_47e56b81_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_30e129c3_result_delayed_u0<=1'h0;
else reg_30e129c3_result_delayed_u0<=reg_30e129c3_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_46b7b9ba_result_delayed_u0<=1'h0;
else reg_46b7b9ba_result_delayed_u0<=reg_46b7b9ba_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_005750dc_result_delayed_result_delayed_u0<=1'h0;
else reg_005750dc_result_delayed_result_delayed_u0<=reg_005750dc_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5236af83_result_delayed_u0<=1'h0;
else reg_5236af83_result_delayed_u0<=reg_5236af83_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_029c8613_result_delayed_result_delayed_u0<=1'h0;
else reg_029c8613_result_delayed_result_delayed_u0<=reg_029c8613_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_69b415a1_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_69b415a1_result_delayed_result_delayed_result_delayed_u0<=reg_69b415a1_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6a850ff6_result_delayed_u0<=1'h0;
else reg_6a850ff6_result_delayed_u0<=reg_6a850ff6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1f3d20af_u0<=1'h0;
else reg_1f3d20af_u0<=reg_12e4f0a0_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4ef81ecb_result_delayed_u0<=1'h0;
else reg_4ef81ecb_result_delayed_u0<=reg_4ef81ecb_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a5ce622_result_delayed_u0<=1'h0;
else reg_7a5ce622_result_delayed_u0<=reg_7a5ce622_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6efe4388_result_delayed_result_delayed_u0<=1'h0;
else reg_6efe4388_result_delayed_result_delayed_u0<=reg_6efe4388_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7b991f92_result_delayed_result_delayed_u0<=1'h0;
else reg_7b991f92_result_delayed_result_delayed_u0<=reg_7b991f92_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_12bc27dd_result_delayed_result_delayed_u0<=1'h0;
else reg_12bc27dd_result_delayed_result_delayed_u0<=reg_12bc27dd_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4bc316c8_result_delayed_u0<=1'h0;
else reg_4bc316c8_result_delayed_u0<=reg_4bc316c8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_33a8b808_u0<=1'h0;
else reg_33a8b808_u0<=reg_19b1e534_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_63cbe06a_u0<=1'h0;
else reg_63cbe06a_u0<=reg_0bd5de0a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1795d1e7_result_delayed_u0<=1'h0;
else reg_1795d1e7_result_delayed_u0<=reg_1795d1e7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3126cd62_result_delayed_u0<=1'h0;
else reg_3126cd62_result_delayed_u0<=reg_3126cd62_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_37b15a18_result_delayed_result_delayed_u0<=1'h0;
else reg_37b15a18_result_delayed_result_delayed_u0<=reg_37b15a18_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1324a63d_result_delayed_result_delayed_u0<=1'h0;
else reg_1324a63d_result_delayed_result_delayed_u0<=reg_1324a63d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3db3d453_result_delayed_u0<=1'h0;
else reg_3db3d453_result_delayed_u0<=reg_3db3d453_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_697bf970_result_delayed_u0<=1'h0;
else reg_697bf970_result_delayed_u0<=reg_697bf970_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_51cd934d_result_delayed_u0<=1'h0;
else reg_51cd934d_result_delayed_u0<=reg_51cd934d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1554b782_result_delayed_result_delayed_u0<=1'h0;
else reg_1554b782_result_delayed_result_delayed_u0<=reg_1554b782_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0f0fdd38_result_delayed_u0<=1'h0;
else reg_0f0fdd38_result_delayed_u0<=reg_0f0fdd38_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_45a71573_result_delayed_u0<=1'h0;
else reg_45a71573_result_delayed_u0<=reg_45a71573_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_12e4f0a0_result_delayed_u0<=1'h0;
else reg_12e4f0a0_result_delayed_u0<=reg_12e4f0a0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_34478ce7_result_delayed_u0<=1'h0;
else reg_34478ce7_result_delayed_u0<=reg_34478ce7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3b9cf399_result_delayed_u0<=1'h0;
else reg_3b9cf399_result_delayed_u0<=reg_3b9cf399_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1ec2c3a2_result_delayed_u0<=1'h0;
else reg_1ec2c3a2_result_delayed_u0<=reg_1ec2c3a2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4fad7ce4_result_delayed_u0<=1'h0;
else reg_4fad7ce4_result_delayed_u0<=reg_4fad7ce4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_16e37f2c_result_delayed_u0<=1'h0;
else reg_16e37f2c_result_delayed_u0<=reg_16e37f2c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_25cb699d_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_25cb699d_result_delayed_result_delayed_result_delayed_u0<=reg_25cb699d_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_19b1e534_result_delayed_u0<=1'h0;
else reg_19b1e534_result_delayed_u0<=reg_19b1e534_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_787cb445_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_787cb445_result_delayed_result_delayed_result_delayed_u0<=reg_787cb445_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6768af3f_result_delayed_u0<=1'h0;
else reg_6768af3f_result_delayed_u0<=reg_6768af3f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7d7ca566_result_delayed_u0<=1'h0;
else reg_7d7ca566_result_delayed_u0<=reg_7d7ca566_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_65dbefa4_result_delayed_u0<=1'h0;
else reg_65dbefa4_result_delayed_u0<=reg_65dbefa4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0924240b_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_0924240b_result_delayed_result_delayed_result_delayed_u0<=reg_0924240b_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_40f3fed8_result_delayed_u0<=1'h0;
else reg_40f3fed8_result_delayed_u0<=reg_40f3fed8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0f03e5b9_result_delayed_u0<=1'h0;
else reg_0f03e5b9_result_delayed_u0<=reg_0f03e5b9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7cb11462_result_delayed_result_delayed_u0<=1'h0;
else reg_7cb11462_result_delayed_result_delayed_u0<=reg_7cb11462_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_29f9ddea_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_29f9ddea_result_delayed_result_delayed_result_delayed_u0<=reg_29f9ddea_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2bd5f75e_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_2bd5f75e_result_delayed_result_delayed_result_delayed_u0<=reg_2bd5f75e_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_52798be3_result_delayed_u0<=1'h0;
else reg_52798be3_result_delayed_u0<=reg_52798be3_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_09f461a1_result_delayed_result_delayed_u0<=1'h0;
else reg_09f461a1_result_delayed_result_delayed_u0<=reg_09f461a1_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_633a5b40_result_delayed_u0<=1'h0;
else reg_633a5b40_result_delayed_u0<=reg_633a5b40_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1ba0d353_result_delayed_u0<=1'h0;
else reg_1ba0d353_result_delayed_u0<=reg_1ba0d353_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7b9f9b79_result_delayed_u0<=1'h0;
else reg_7b9f9b79_result_delayed_u0<=reg_7b9f9b79_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_10d31157_result_delayed_u0<=1'h0;
else reg_10d31157_result_delayed_u0<=reg_10d31157_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_368fce58_result_delayed_u0<=1'h0;
else reg_368fce58_result_delayed_u0<=reg_368fce58_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2ae45e03_result_delayed_result_delayed_u0<=1'h0;
else reg_2ae45e03_result_delayed_result_delayed_u0<=reg_2ae45e03_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_79ff2594_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_79ff2594_result_delayed_result_delayed_result_delayed_u0<=reg_79ff2594_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_12299b2b_result_delayed_u0<=1'h0;
else reg_12299b2b_result_delayed_u0<=reg_12299b2b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0bd5de0a_result_delayed_u0<=1'h0;
else reg_0bd5de0a_result_delayed_u0<=reg_0bd5de0a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_32d59a7c_result_delayed_u0<=1'h0;
else reg_32d59a7c_result_delayed_u0<=reg_32d59a7c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7834905a_result_delayed_u0<=1'h0;
else reg_7834905a_result_delayed_u0<=reg_7834905a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_039f5f0f_result_delayed_u0<=1'h0;
else reg_039f5f0f_result_delayed_u0<=reg_039f5f0f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_04a958f3_result_delayed_result_delayed_u0<=1'h0;
else reg_04a958f3_result_delayed_result_delayed_u0<=reg_04a958f3_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4ef81ecb_result_delayed_result_delayed_u0<=1'h0;
else reg_4ef81ecb_result_delayed_result_delayed_u0<=reg_4ef81ecb_result_delayed_u0;
end
assign or_u1106_u0=and_u3611_u0|and_u3610_u0;
assign mux_u360=(and_u3611_u0)?1'h1:1'h0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_787cb445_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_787cb445_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_787cb445_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1801415e_result_delayed_result_delayed_u0<=1'h0;
else reg_1801415e_result_delayed_result_delayed_u0<=reg_1801415e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_11cd6f36_result_delayed_u0<=1'h0;
else reg_11cd6f36_result_delayed_u0<=reg_11cd6f36_u0;
end
assign mux_u361_u0=(and_u3614_u0)?1'h1:mux_u360;
assign or_u1107_u0=and_u3614_u0|or_u1106_u0;
assign or_u1108_u0=and_u3614_u0|and_u3611_u0;
assign mux_u362_u0=(and_u3614_u0)?32'h4:32'h200;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4e481e21_u0<=1'h0;
else reg_4e481e21_u0<=reg_3a07cc10_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2258ca11_u0<=1'h0;
else reg_2258ca11_u0<=reg_4e481e21_result_delayed_result_delayed_u0;
end
assign or_u1109_u0=and_u3614_u0|and_u3611_u0;
assign and_u3613_u0=and_u3605_u0&and_u3616_u0;
assign or_u1110_u0=reg_2258ca11_u0|or_u1105_u0;
assign or_u1111_u0=and_u3614_u0|and_u3611_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4e481e21_result_delayed_u0<=1'h0;
else reg_4e481e21_result_delayed_u0<=reg_4e481e21_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3a07cc10_u0<=1'h0;
else reg_3a07cc10_u0<=and_u3614_u0;
end
assign or_u1112_u0=and_u3614_u0|and_u3611_u0;
assign and_u3614_u0=and_u3604_u0&and_u3616_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4e481e21_result_delayed_result_delayed_u0<=1'h0;
else reg_4e481e21_result_delayed_result_delayed_u0<=reg_4e481e21_result_delayed_u0;
end
assign and_u3615_u0=and_u3603_u0&and_u3634_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u240_u0<=1'h0;
else and_delayed_u240_u0<=and_u3615_u0;
end
assign or_u1113_u0=or_u1110_u0|and_delayed_u240_u0;
assign and_u3616_u0=and_u3602_u0&and_u3634_u0;
assign equals_u190_a_signed={31'b0, port_5b3d11e3_};
assign equals_u190_b_signed=32'h1;
assign equals_u190=equals_u190_a_signed==equals_u190_b_signed;
assign and_u3617_u0=and_u3634_u0&equals_u190;
assign not_u590_u0=~equals_u190;
assign and_u3618_u0=and_u3634_u0&not_u590_u0;
assign and_u3619_u0=and_u3633_u0&port_02986e5e_;
assign not_u591_u0=~port_02986e5e_;
assign and_u3620_u0=and_u3633_u0&not_u591_u0;
assign lessThan_u87_a_signed=port_5aad7090_;
assign lessThan_u87_b_signed=port_598dd3c9_;
assign lessThan_u87=lessThan_u87_a_signed<lessThan_u87_b_signed;
assign not_u592_u0=~lessThan_u87;
assign and_u3621_u0=and_u3630_u0&lessThan_u87;
assign and_u3622_u0=and_u3630_u0&not_u592_u0;
assign and_u3623_u0=and_u3628_u0&not_u593_u0;
assign not_u593_u0=~port_19d5fffb_;
assign and_u3624_u0=and_u3628_u0&port_19d5fffb_;
assign add=port_5aad7090_+32'h0;
assign and_u3625_u0=and_u3626_u0&port_680d32a7_;
assign simplePinWrite_u518=and_u3626_u0&{1{and_u3626_u0}};
assign simplePinWrite_u519=16'h1&{16{1'h1}};
assign simplePinWrite_u520=port_7e2c6053_;
assign add_u476=port_5aad7090_+32'h1;
always @(posedge CLK)
begin
if (and_u3626_u0)
syncEnable_u688<=port_7e2c6053_;
end
assign and_u3626_u0=and_u3624_u0&and_u3628_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u241_u0<=1'h0;
else and_delayed_u241_u0<=and_u3626_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_22db32bc_u0<=1'h0;
else reg_22db32bc_u0<=and_u3627_u0;
end
assign and_u3627_u0=and_u3623_u0&and_u3628_u0;
assign mux_u363_u0=(reg_22db32bc_u0)?syncEnable_u689_u0:syncEnable_u688;
always @(posedge CLK)
begin
if (and_u3628_u0)
syncEnable_u689_u0<=mux_u375_u0;
end
assign and_u3628_u0=and_u3621_u0&and_u3630_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u242_u0<=1'h0;
else and_delayed_u242_u0<=and_u3628_u0;
end
assign mux_u364_u0=(and_delayed_u243_u0)?syncEnable_u690_u0:mux_u363_u0;
assign and_u3629_u0=and_u3622_u0&and_u3630_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u243_u0<=1'h0;
else and_delayed_u243_u0<=and_u3629_u0;
end
assign mux_u365_u0=(and_delayed_u243_u0)?32'h0:syncEnable_u691_u0;
always @(posedge CLK)
begin
if (and_u3630_u0)
syncEnable_u690_u0<=mux_u375_u0;
end
always @(posedge CLK)
begin
if (and_u3630_u0)
syncEnable_u691_u0<=mux_u374_u0;
end
assign mux_u366_u0=(and_delayed_u244_u0)?mux_u365_u0:syncEnable_u692_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_10a5074b_u0<=1'h0;
else reg_10a5074b_u0<=and_u3631_u0;
end
assign mux_u367_u0=(and_delayed_u244_u0)?mux_u364_u0:syncEnable_u693_u0;
always @(posedge CLK)
begin
if (and_u3633_u0)
syncEnable_u692_u0<=mux_u374_u0;
end
assign and_u3630_u0=and_u3619_u0&and_u3633_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u244_u0<=1'h0;
else and_delayed_u244_u0<=and_u3630_u0;
end
always @(posedge CLK)
begin
if (and_u3633_u0)
syncEnable_u693_u0<=mux_u375_u0;
end
assign and_u3631_u0=and_u3620_u0&and_u3633_u0;
always @(posedge CLK)
begin
if (and_u3634_u0)
syncEnable_u694_u0<=mux_u375_u0;
end
assign and_u3632_u0=and_u3618_u0&and_u3634_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u245_u0<=1'h0;
else and_delayed_u245_u0<=and_u3632_u0;
end
assign and_u3633_u0=and_u3617_u0&and_u3634_u0;
assign mux_u368_u0=(and_delayed_u245_u0)?syncEnable_u695_u0:mux_u366_u0;
always @(posedge CLK)
begin
if (and_u3634_u0)
syncEnable_u695_u0<=mux_u374_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u246_u0<=1'h0;
else and_delayed_u246_u0<=and_u3633_u0;
end
assign mux_u369_u0=(and_delayed_u245_u0)?syncEnable_u694_u0:mux_u367_u0;
assign mux_u370_u0=(or_u1109_u0)?32'h0:add_u476;
assign or_u1114_u0=or_u1109_u0|and_u3626_u0;
assign latch_512b7f83_out=(block_GO_delayed_u12)?mux_u368_u0:latch_512b7f83_reg;
always @(posedge CLK)
begin
if (block_GO_delayed_u12)
latch_512b7f83_reg<=mux_u368_u0;
end
always @(posedge CLK)
begin
if (block_GO_delayed_u12)
latch_57dc3c15_reg<=mux_u369_u0;
end
assign latch_57dc3c15_out=(block_GO_delayed_u12)?mux_u369_u0:latch_57dc3c15_reg;
assign or_u1115_u0=or_u1107_u0|and_u3629_u0;
assign mux_u371_u0=(or_u1107_u0)?mux_u361_u0:1'h0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
block_GO_delayed_u12<=1'h0;
else block_GO_delayed_u12<=and_u3634_u0;
end
assign mux_u372_u0=(or_u1108_u0)?{22'b0, mux_u362_u0[9], 6'b0, mux_u362_u0[2], 2'b0}:32'hffffffff;
assign or_u1116_u0=or_u1108_u0|and_u3629_u0;
assign or_u1117_u0=or_u1112_u0|and_u3629_u0;
assign mux_u373_u0=(or_u1112_u0)?1'h1:1'h0;
assign and_u3634_u0=or_u1118_u0&or_u1118_u0;
always @(posedge CLK or posedge syncEnable_u696_u0)
begin
if (syncEnable_u696_u0)
loopControl_u9<=1'h0;
else loopControl_u9<=or_u1113_u0;
end
assign or_u1118_u0=loopControl_u9|reg_7a06e94d_result_delayed_u0;
always @(posedge CLK)
begin
if (reg_7a06e94d_result_delayed_u0)
syncEnable_u696_u0<=RESET;
end
always @(posedge CLK)
begin
if (or_u1113_u0)
fbReg_Out1Portvalue_u4<=latch_57dc3c15_out;
end
always @(posedge CLK)
begin
if (or_u1113_u0)
fbReg_temp_fsmOldState_resized_LH2_xy_7_u0<=latch_512b7f83_out;
end
assign mux_u374_u0=(loopControl_u9)?fbReg_temp_fsmOldState_resized_LH2_xy_7_u0:32'h0;
assign mux_u375_u0=(loopControl_u9)?fbReg_Out1Portvalue_u4:16'h0;
assign or_u1119_u0=GO|or_u1117_u0;
assign mux_u376_u0=(GO)?1'h0:mux_u373_u0;
assign mux_u377_u0=(GO)?1'h0:mux_u371_u0;
assign or_u1120_u0=GO|or_u1115_u0;
assign or_u1121_u0=GO|or_u1111_u0;
assign or_u1122_u0=GO|or_u1114_u0;
assign mux_u378_u0=(GO)?32'h0:mux_u370_u0;
assign mux_u379_u0=(GO)?32'hffffffff:mux_u372_u0;
assign or_u1123_u0=GO|or_u1116_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a06e94d_u0<=1'h0;
else reg_7a06e94d_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a06e94d_result_delayed_u0<=1'h0;
else reg_7a06e94d_result_delayed_u0<=reg_7a06e94d_u0;
end
assign RESULT=or_u1121_u0;
assign RESULT_u2119=32'h0;
assign RESULT_u2120=or_u1120_u0;
assign RESULT_u2121=mux_u377_u0;
assign RESULT_u2122=or_u1122_u0;
assign RESULT_u2123=mux_u378_u0;
assign RESULT_u2124=or_u1123_u0;
assign RESULT_u2125=mux_u379_u0;
assign RESULT_u2126=or_u1119_u0;
assign RESULT_u2127=mux_u376_u0;
assign RESULT_u2128=and_u3626_u0;
assign RESULT_u2129=add;
assign RESULT_u2130=3'h1;
assign RESULT_u2131=simplePinWrite_u518;
assign RESULT_u2132=simplePinWrite_u519;
assign RESULT_u2133=simplePinWrite_u516;
assign RESULT_u2134=simplePinWrite;
assign RESULT_u2135=simplePinWrite_u517;
assign RESULT_u2136=simplePinWrite_u520;
assign DONE=1'h0;
endmodule



module resized_LH2_xy_endianswapper_4f771850_(endianswapper_4f771850_in, endianswapper_4f771850_out);
input	[15:0]	endianswapper_4f771850_in;
output	[15:0]	endianswapper_4f771850_out;
assign endianswapper_4f771850_out=endianswapper_4f771850_in;
endmodule



module resized_LH2_xy_endianswapper_11152082_(endianswapper_11152082_in, endianswapper_11152082_out);
input	[15:0]	endianswapper_11152082_in;
output	[15:0]	endianswapper_11152082_out;
assign endianswapper_11152082_out=endianswapper_11152082_in;
endmodule



module resized_LH2_xy_stateVar_rowRepeated(bus_2fffcdc9_, bus_1df4e7c6_, bus_543e42b8_, bus_3f0e41dd_, bus_558d89ec_, bus_6faa67c2_, bus_45cec17e_);
input		bus_2fffcdc9_;
input		bus_1df4e7c6_;
input		bus_543e42b8_;
input	[15:0]	bus_3f0e41dd_;
input		bus_558d89ec_;
input	[15:0]	bus_6faa67c2_;
output	[15:0]	bus_45cec17e_;
wire		or_0ecb9eec_u0;
wire	[15:0]	endianswapper_4f771850_out;
wire	[15:0]	endianswapper_11152082_out;
reg	[15:0]	stateVar_rowRepeated_u4=16'h1;
wire	[15:0]	mux_7e53af3d_u0;
assign or_0ecb9eec_u0=bus_543e42b8_|bus_558d89ec_;
resized_LH2_xy_endianswapper_4f771850_ resized_LH2_xy_endianswapper_4f771850__1(.endianswapper_4f771850_in(mux_7e53af3d_u0), 
  .endianswapper_4f771850_out(endianswapper_4f771850_out));
resized_LH2_xy_endianswapper_11152082_ resized_LH2_xy_endianswapper_11152082__1(.endianswapper_11152082_in(stateVar_rowRepeated_u4), 
  .endianswapper_11152082_out(endianswapper_11152082_out));
assign bus_45cec17e_=endianswapper_11152082_out;
always @(posedge bus_2fffcdc9_ or posedge bus_1df4e7c6_)
begin
if (bus_1df4e7c6_)
stateVar_rowRepeated_u4<=16'h1;
else if (or_0ecb9eec_u0)
stateVar_rowRepeated_u4<=endianswapper_4f771850_out;
end
assign mux_7e53af3d_u0=(bus_543e42b8_)?bus_3f0e41dd_:16'h1;
endmodule



module resized_LH2_xy_forge_memory_512x16_38(CLK, EN, WE, ADDR, DIN, DOUT, DONE);
input		CLK;
input		EN;
input		WE;
input	[31:0]	ADDR;
input	[15:0]	DIN;
output	[15:0]	DOUT;
output		DONE;
wire		we_0;
wire	[15:0]	pre_dout_0;
wire		we_1;
wire	[15:0]	pre_dout_1;
wire		we_2;
wire	[15:0]	pre_dout_2;
wire		we_3;
wire	[15:0]	pre_dout_3;
reg	[15:0]	mux_out;
reg		wen_done;
assign we_0=WE&(ADDR[31:7]==25'h0);
assign we_1=WE&(ADDR[31:7]==25'h1);
assign we_2=WE&(ADDR[31:7]==25'h2);
assign we_3=WE&(ADDR[31:7]==25'h3);
always @(ADDR or pre_dout_0 or pre_dout_1 or pre_dout_2 or pre_dout_3)
begin
case (ADDR[31:7])25'd0:mux_out=pre_dout_0;
25'd1:mux_out=pre_dout_1;
25'd2:mux_out=pre_dout_2;
25'd3:mux_out=pre_dout_3;
default:mux_out=16'h0;
endcase end
always @(posedge CLK)
begin
wen_done<=WE;
end
assign DOUT=mux_out;
assign DONE=EN&!WE|wen_done;
//  Memory array element: COL: 0, ROW: 0
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_256(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[0]), .O(pre_dout_0[0]));
//  Memory array element: COL: 0, ROW: 1
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_257(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[1]), .O(pre_dout_0[1]));
//  Memory array element: COL: 0, ROW: 2
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_258(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[2]), .O(pre_dout_0[2]));
//  Memory array element: COL: 0, ROW: 3
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_259(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[3]), .O(pre_dout_0[3]));
//  Memory array element: COL: 0, ROW: 4
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_260(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[4]), .O(pre_dout_0[4]));
//  Memory array element: COL: 0, ROW: 5
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_261(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[5]), .O(pre_dout_0[5]));
//  Memory array element: COL: 0, ROW: 6
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_262(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[6]), .O(pre_dout_0[6]));
//  Memory array element: COL: 0, ROW: 7
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_263(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[7]), .O(pre_dout_0[7]));
//  Memory array element: COL: 0, ROW: 8
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_264(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[8]), .O(pre_dout_0[8]));
//  Memory array element: COL: 0, ROW: 9
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_265(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[9]), .O(pre_dout_0[9]));
//  Memory array element: COL: 0, ROW: 10
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_266(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[10]), .O(pre_dout_0[10]));
//  Memory array element: COL: 0, ROW: 11
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_267(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[11]), .O(pre_dout_0[11]));
//  Memory array element: COL: 0, ROW: 12
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_268(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[12]), .O(pre_dout_0[12]));
//  Memory array element: COL: 0, ROW: 13
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_269(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[13]), .O(pre_dout_0[13]));
//  Memory array element: COL: 0, ROW: 14
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_270(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[14]), .O(pre_dout_0[14]));
//  Memory array element: COL: 0, ROW: 15
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_271(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[15]), .O(pre_dout_0[15]));
//  Memory array element: COL: 1, ROW: 0
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_272(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[0]), .O(pre_dout_1[0]));
//  Memory array element: COL: 1, ROW: 1
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_273(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[1]), .O(pre_dout_1[1]));
//  Memory array element: COL: 1, ROW: 2
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_274(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[2]), .O(pre_dout_1[2]));
//  Memory array element: COL: 1, ROW: 3
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_275(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[3]), .O(pre_dout_1[3]));
//  Memory array element: COL: 1, ROW: 4
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_276(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[4]), .O(pre_dout_1[4]));
//  Memory array element: COL: 1, ROW: 5
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_277(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[5]), .O(pre_dout_1[5]));
//  Memory array element: COL: 1, ROW: 6
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_278(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[6]), .O(pre_dout_1[6]));
//  Memory array element: COL: 1, ROW: 7
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_279(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[7]), .O(pre_dout_1[7]));
//  Memory array element: COL: 1, ROW: 8
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_280(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[8]), .O(pre_dout_1[8]));
//  Memory array element: COL: 1, ROW: 9
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_281(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[9]), .O(pre_dout_1[9]));
//  Memory array element: COL: 1, ROW: 10
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_282(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[10]), .O(pre_dout_1[10]));
//  Memory array element: COL: 1, ROW: 11
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_283(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[11]), .O(pre_dout_1[11]));
//  Memory array element: COL: 1, ROW: 12
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_284(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[12]), .O(pre_dout_1[12]));
//  Memory array element: COL: 1, ROW: 13
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_285(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[13]), .O(pre_dout_1[13]));
//  Memory array element: COL: 1, ROW: 14
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_286(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[14]), .O(pre_dout_1[14]));
//  Memory array element: COL: 1, ROW: 15
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_287(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[15]), .O(pre_dout_1[15]));
//  Memory array element: COL: 2, ROW: 0
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_288(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[0]), .O(pre_dout_2[0]));
//  Memory array element: COL: 2, ROW: 1
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_289(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[1]), .O(pre_dout_2[1]));
//  Memory array element: COL: 2, ROW: 2
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_290(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[2]), .O(pre_dout_2[2]));
//  Memory array element: COL: 2, ROW: 3
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_291(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[3]), .O(pre_dout_2[3]));
//  Memory array element: COL: 2, ROW: 4
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_292(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[4]), .O(pre_dout_2[4]));
//  Memory array element: COL: 2, ROW: 5
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_293(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[5]), .O(pre_dout_2[5]));
//  Memory array element: COL: 2, ROW: 6
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_294(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[6]), .O(pre_dout_2[6]));
//  Memory array element: COL: 2, ROW: 7
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_295(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[7]), .O(pre_dout_2[7]));
//  Memory array element: COL: 2, ROW: 8
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_296(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[8]), .O(pre_dout_2[8]));
//  Memory array element: COL: 2, ROW: 9
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_297(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[9]), .O(pre_dout_2[9]));
//  Memory array element: COL: 2, ROW: 10
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_298(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[10]), .O(pre_dout_2[10]));
//  Memory array element: COL: 2, ROW: 11
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_299(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[11]), .O(pre_dout_2[11]));
//  Memory array element: COL: 2, ROW: 12
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_300(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[12]), .O(pre_dout_2[12]));
//  Memory array element: COL: 2, ROW: 13
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_301(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[13]), .O(pre_dout_2[13]));
//  Memory array element: COL: 2, ROW: 14
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_302(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[14]), .O(pre_dout_2[14]));
//  Memory array element: COL: 2, ROW: 15
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_303(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[15]), .O(pre_dout_2[15]));
//  Memory array element: COL: 3, ROW: 0
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_304(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[0]), .O(pre_dout_3[0]));
//  Memory array element: COL: 3, ROW: 1
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_305(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[1]), .O(pre_dout_3[1]));
//  Memory array element: COL: 3, ROW: 2
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_306(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[2]), .O(pre_dout_3[2]));
//  Memory array element: COL: 3, ROW: 3
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_307(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[3]), .O(pre_dout_3[3]));
//  Memory array element: COL: 3, ROW: 4
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_308(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[4]), .O(pre_dout_3[4]));
//  Memory array element: COL: 3, ROW: 5
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_309(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[5]), .O(pre_dout_3[5]));
//  Memory array element: COL: 3, ROW: 6
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_310(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[6]), .O(pre_dout_3[6]));
//  Memory array element: COL: 3, ROW: 7
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_311(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[7]), .O(pre_dout_3[7]));
//  Memory array element: COL: 3, ROW: 8
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_312(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[8]), .O(pre_dout_3[8]));
//  Memory array element: COL: 3, ROW: 9
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_313(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[9]), .O(pre_dout_3[9]));
//  Memory array element: COL: 3, ROW: 10
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_314(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[10]), .O(pre_dout_3[10]));
//  Memory array element: COL: 3, ROW: 11
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_315(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[11]), .O(pre_dout_3[11]));
//  Memory array element: COL: 3, ROW: 12
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_316(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[12]), .O(pre_dout_3[12]));
//  Memory array element: COL: 3, ROW: 13
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_317(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[13]), .O(pre_dout_3[13]));
//  Memory array element: COL: 3, ROW: 14
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_318(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[14]), .O(pre_dout_3[14]));
//  Memory array element: COL: 3, ROW: 15
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_319(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[15]), .O(pre_dout_3[15]));
endmodule



module resized_LH2_xy_structuralmemory_10a0b0c5_(CLK_u20, bus_5a27453b_, bus_2abe7aae_, bus_3da3e1e4_, bus_0a872caa_, bus_4328a1e0_, bus_12b5a8c1_, bus_2b80c1a2_, bus_2bfcb357_);
input		CLK_u20;
input		bus_5a27453b_;
input	[31:0]	bus_2abe7aae_;
input	[2:0]	bus_3da3e1e4_;
input		bus_0a872caa_;
input		bus_4328a1e0_;
input	[15:0]	bus_12b5a8c1_;
output	[15:0]	bus_2b80c1a2_;
output		bus_2bfcb357_;
wire		or_58a44447_u0;
wire	[15:0]	bus_1827f4c7_;
wire		or_5c9e58f4_u0;
wire		not_344a32a6_u0;
wire		and_351ffe6d_u0;
reg		logicalMem_123f0e02_we_delay0_u0=1'h0;
assign or_58a44447_u0=bus_0a872caa_|bus_4328a1e0_;
resized_LH2_xy_forge_memory_512x16_38 resized_LH2_xy_forge_memory_512x16_38_instance0(.CLK(CLK_u20), 
  .EN(or_58a44447_u0), .WE(bus_4328a1e0_), .ADDR(bus_2abe7aae_), .DIN(bus_12b5a8c1_), 
  .DOUT(bus_1827f4c7_), .DONE());
assign or_5c9e58f4_u0=and_351ffe6d_u0|logicalMem_123f0e02_we_delay0_u0;
assign not_344a32a6_u0=~bus_4328a1e0_;
assign bus_2b80c1a2_=bus_1827f4c7_;
assign bus_2bfcb357_=or_5c9e58f4_u0;
assign and_351ffe6d_u0=bus_0a872caa_&not_344a32a6_u0;
always @(posedge CLK_u20 or posedge bus_5a27453b_)
begin
if (bus_5a27453b_)
logicalMem_123f0e02_we_delay0_u0<=1'h0;
else logicalMem_123f0e02_we_delay0_u0<=bus_4328a1e0_;
end
endmodule



module resized_LH2_xy_reset(CLK, RESET, GO, RESULT, RESULT_u2137, RESULT_u2138, RESULT_u2139, DONE);
input		CLK;
input		RESET;
input		GO;
output		RESULT;
output	[15:0]	RESULT_u2137;
output		RESULT_u2138;
output	[15:0]	RESULT_u2139;
output		DONE;
reg		reg_468aabc3_u0=1'h0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_468aabc3_u0<=1'h0;
else reg_468aabc3_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u2137=16'h1;
assign RESULT_u2138=GO;
assign RESULT_u2139=16'h0;
assign DONE=reg_468aabc3_u0;
endmodule



module resized_LH2_xy_globalreset_physical_0b41fdb2_(bus_0a890099_, bus_132690ba_, bus_112f0657_);
input		bus_0a890099_;
input		bus_132690ba_;
output		bus_112f0657_;
reg		cross_u41=1'h0;
wire		not_15889bba_u0;
reg		final_u41=1'h1;
reg		glitch_u41=1'h0;
wire		or_01bf3353_u0;
reg		sample_u41=1'h0;
wire		and_7e7040bf_u0;
always @(posedge bus_0a890099_)
begin
cross_u41<=sample_u41;
end
assign not_15889bba_u0=~and_7e7040bf_u0;
assign bus_112f0657_=or_01bf3353_u0;
always @(posedge bus_0a890099_)
begin
final_u41<=not_15889bba_u0;
end
always @(posedge bus_0a890099_)
begin
glitch_u41<=cross_u41;
end
assign or_01bf3353_u0=bus_132690ba_|final_u41;
always @(posedge bus_0a890099_)
begin
sample_u41<=1'h1;
end
assign and_7e7040bf_u0=cross_u41&glitch_u41;
endmodule



module resized_LH2_xy_consumeRow(CLK, RESET, GO, port_174a8800_, port_19cd6551_, port_29086a48_, port_21dccef2_, RESULT, RESULT_u2140, RESULT_u2141, RESULT_u2142, RESULT_u2143, RESULT_u2144, RESULT_u2145, RESULT_u2146, RESULT_u2147, RESULT_u2148, RESULT_u2149, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_174a8800_;
input		port_19cd6551_;
input		port_29086a48_;
input	[15:0]	port_21dccef2_;
output		RESULT;
output	[15:0]	RESULT_u2140;
output		RESULT_u2141;
output	[31:0]	RESULT_u2142;
output	[15:0]	RESULT_u2143;
output	[2:0]	RESULT_u2144;
output		RESULT_u2145;
output	[31:0]	RESULT_u2146;
output	[15:0]	RESULT_u2147;
output	[2:0]	RESULT_u2148;
output		RESULT_u2149;
output		DONE;
wire		simplePinWrite;
wire	[31:0]	add;
wire	[31:0]	add_u477;
reg		reg_7939cf59_u0=1'h0;
wire		or_u1124_u0;
wire		and_u3635_u0;
wire	[15:0]	add_u478;
reg	[15:0]	syncEnable_u697=16'h0;
reg		reg_5f4f6df8_u0=1'h0;
wire		and_u3636_u0;
wire		lessThanEqualTo;
wire signed	[16:0]	lessThanEqualTo_a_signed;
wire signed	[16:0]	lessThanEqualTo_b_signed;
wire		not_u594_u0;
wire		and_u3637_u0;
wire		and_u3638_u0;
wire		and_u3639_u0;
wire	[15:0]	latch_02831c6f_out;
reg	[15:0]	latch_02831c6f_reg=16'h0;
wire	[15:0]	mux_u380;
wire		or_u1125_u0;
wire	[15:0]	add_u479;
wire		and_u3640_u0;
wire		and_u3641_u0;
wire		lessThanEqualTo_u4;
wire signed	[16:0]	lessThanEqualTo_u4_b_signed;
wire signed	[16:0]	lessThanEqualTo_u4_a_signed;
wire		and_u3642_u0;
wire		not_u595_u0;
wire		and_u3643_u0;
reg		and_delayed_u247=1'h0;
wire	[15:0]	subtract;
wire	[31:0]	add_u480;
wire		or_u1126_u0;
reg		reg_0b1bb952_u0=1'h0;
wire		and_u3644_u0;
wire	[15:0]	add_u481;
reg	[15:0]	syncEnable_u698_u0=16'h0;
wire		or_u1127_u0;
reg	[15:0]	latch_301cd5cd_reg=16'h0;
wire	[15:0]	latch_301cd5cd_out;
wire	[15:0]	mux_u381_u0;
reg	[15:0]	syncEnable_u699_u0=16'h0;
reg		reg_307b44a0_u0=1'h0;
assign simplePinWrite=GO&{1{GO}};
assign add={14'b0, port_174a8800_, 2'b0}+{mux_u380[15], mux_u380[15], mux_u380[15], mux_u380[15], mux_u380[15], mux_u380[15], mux_u380[15], mux_u380[15], mux_u380[15], mux_u380[15], mux_u380[15], mux_u380[15], mux_u380[15], mux_u380[15], mux_u380[15], mux_u380[15], mux_u380};
assign add_u477={add[19], add[19], add[19], add[19], add[19], add[19], add[19], add[19], add[19], add[19], add[19], add[19], add[19:0]}+32'h0;
always @(posedge CLK or posedge and_u3636_u0 or posedge or_u1124_u0)
begin
if (or_u1124_u0)
reg_7939cf59_u0<=1'h0;
else if (and_u3636_u0)
reg_7939cf59_u0<=1'h1;
else reg_7939cf59_u0<=reg_7939cf59_u0;
end
assign or_u1124_u0=and_u3635_u0|RESET;
assign and_u3635_u0=reg_7939cf59_u0&port_29086a48_;
assign add_u478=mux_u380+16'h1;
always @(posedge CLK)
begin
if (and_u3636_u0)
syncEnable_u697<=add_u478;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5f4f6df8_u0<=1'h0;
else reg_5f4f6df8_u0<=and_u3636_u0;
end
assign and_u3636_u0=and_u3638_u0&or_u1125_u0;
assign lessThanEqualTo_a_signed={mux_u380[15], mux_u380};
assign lessThanEqualTo_b_signed=17'h3;
assign lessThanEqualTo=lessThanEqualTo_a_signed<=lessThanEqualTo_b_signed;
assign not_u594_u0=~lessThanEqualTo;
assign and_u3637_u0=or_u1125_u0&not_u594_u0;
assign and_u3638_u0=or_u1125_u0&lessThanEqualTo;
assign and_u3639_u0=and_u3637_u0&or_u1125_u0;
assign latch_02831c6f_out=(GO)?port_21dccef2_:latch_02831c6f_reg;
always @(posedge CLK)
begin
if (GO)
latch_02831c6f_reg<=port_21dccef2_;
end
assign mux_u380=(reg_5f4f6df8_u0)?syncEnable_u697:16'h0;
assign or_u1125_u0=reg_5f4f6df8_u0|GO;
assign add_u479=port_174a8800_+16'h1;
assign and_u3640_u0=and_u3642_u0&or_u1127_u0;
assign and_u3641_u0=and_u3643_u0&or_u1127_u0;
assign lessThanEqualTo_u4_a_signed={mux_u381_u0[15], mux_u381_u0};
assign lessThanEqualTo_u4_b_signed=17'h4;
assign lessThanEqualTo_u4=lessThanEqualTo_u4_a_signed<=lessThanEqualTo_u4_b_signed;
assign and_u3642_u0=or_u1127_u0&not_u595_u0;
assign not_u595_u0=~lessThanEqualTo_u4;
assign and_u3643_u0=or_u1127_u0&lessThanEqualTo_u4;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u247<=1'h0;
else and_delayed_u247<=and_u3641_u0;
end
assign subtract=mux_u381_u0-16'h1;
assign add_u480={subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract}+32'h0;
assign or_u1126_u0=and_u3644_u0|RESET;
always @(posedge CLK or posedge and_u3641_u0 or posedge or_u1126_u0)
begin
if (or_u1126_u0)
reg_0b1bb952_u0<=1'h0;
else if (and_u3641_u0)
reg_0b1bb952_u0<=1'h1;
else reg_0b1bb952_u0<=reg_0b1bb952_u0;
end
assign and_u3644_u0=reg_0b1bb952_u0&port_19cd6551_;
assign add_u481=mux_u381_u0+16'h1;
always @(posedge CLK)
begin
if (and_u3641_u0)
syncEnable_u698_u0<=add_u481;
end
assign or_u1127_u0=and_delayed_u247|GO;
always @(posedge CLK)
begin
if (GO)
latch_301cd5cd_reg<=port_21dccef2_;
end
assign latch_301cd5cd_out=(GO)?port_21dccef2_:latch_301cd5cd_reg;
assign mux_u381_u0=(and_delayed_u247)?syncEnable_u698_u0:16'h1;
always @(posedge CLK)
begin
if (GO)
syncEnable_u699_u0<=add_u479;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_307b44a0_u0<=1'h0;
else reg_307b44a0_u0<=and_u3639_u0;
end
assign RESULT=and_u3639_u0;
assign RESULT_u2140=syncEnable_u699_u0;
assign RESULT_u2141=and_u3641_u0;
assign RESULT_u2142=add_u480;
assign RESULT_u2143=latch_301cd5cd_out;
assign RESULT_u2144=3'h1;
assign RESULT_u2145=and_u3636_u0;
assign RESULT_u2146=add_u477;
assign RESULT_u2147=latch_02831c6f_out;
assign RESULT_u2148=3'h1;
assign RESULT_u2149=simplePinWrite;
assign DONE=reg_307b44a0_u0;
endmodule



module resized_LH2_xy_endianswapper_23874674_(endianswapper_23874674_in, endianswapper_23874674_out);
input		endianswapper_23874674_in;
output		endianswapper_23874674_out;
assign endianswapper_23874674_out=endianswapper_23874674_in;
endmodule



module resized_LH2_xy_endianswapper_38de9ae8_(endianswapper_38de9ae8_in, endianswapper_38de9ae8_out);
input		endianswapper_38de9ae8_in;
output		endianswapper_38de9ae8_out;
assign endianswapper_38de9ae8_out=endianswapper_38de9ae8_in;
endmodule



module resized_LH2_xy_stateVar_fsmState_resized_LH2_xy(bus_5fb95275_, bus_4d57ece6_, bus_215b8d1b_, bus_46a6a319_, bus_2a450b51_);
input		bus_5fb95275_;
input		bus_4d57ece6_;
input		bus_215b8d1b_;
input		bus_46a6a319_;
output		bus_2a450b51_;
reg		stateVar_fsmState_resized_LH2_xy_u0=1'h0;
wire		endianswapper_23874674_out;
wire		endianswapper_38de9ae8_out;
always @(posedge bus_5fb95275_ or posedge bus_4d57ece6_)
begin
if (bus_4d57ece6_)
stateVar_fsmState_resized_LH2_xy_u0<=1'h0;
else if (bus_215b8d1b_)
stateVar_fsmState_resized_LH2_xy_u0<=endianswapper_23874674_out;
end
resized_LH2_xy_endianswapper_23874674_ resized_LH2_xy_endianswapper_23874674__1(.endianswapper_23874674_in(bus_46a6a319_), 
  .endianswapper_23874674_out(endianswapper_23874674_out));
resized_LH2_xy_endianswapper_38de9ae8_ resized_LH2_xy_endianswapper_38de9ae8__1(.endianswapper_38de9ae8_in(stateVar_fsmState_resized_LH2_xy_u0), 
  .endianswapper_38de9ae8_out(endianswapper_38de9ae8_out));
assign bus_2a450b51_=endianswapper_38de9ae8_out;
endmodule



module resized_LH2_xy_structuralmemory_57a3ce5d_(CLK_u21, bus_0916e569_, bus_680f5707_, bus_21a49687_, bus_0aab59c9_, bus_3650d95d_, bus_1e93c313_, bus_0f871660_, bus_55b75661_);
input		CLK_u21;
input		bus_0916e569_;
input	[31:0]	bus_680f5707_;
input	[2:0]	bus_21a49687_;
input		bus_0aab59c9_;
input		bus_3650d95d_;
input	[15:0]	bus_1e93c313_;
output	[15:0]	bus_0f871660_;
output		bus_55b75661_;
wire		or_67e4b328_u0;
wire		not_4794121a_u0;
reg		logicalMem_d0e13e1_we_delay0_u0=1'h0;
wire	[15:0]	bus_305dcfd3_;
wire		or_70dee808_u0;
wire		and_635d9962_u0;
assign or_67e4b328_u0=bus_0aab59c9_|bus_3650d95d_;
assign not_4794121a_u0=~bus_3650d95d_;
assign bus_0f871660_=bus_305dcfd3_;
assign bus_55b75661_=or_70dee808_u0;
always @(posedge CLK_u21 or posedge bus_0916e569_)
begin
if (bus_0916e569_)
logicalMem_d0e13e1_we_delay0_u0<=1'h0;
else logicalMem_d0e13e1_we_delay0_u0<=bus_3650d95d_;
end
resized_LH2_xy_forge_memory_512x16_38 resized_LH2_xy_forge_memory_512x16_38_instance1(.CLK(CLK_u21), 
  .EN(or_67e4b328_u0), .WE(bus_3650d95d_), .ADDR(bus_680f5707_), .DIN(bus_1e93c313_), 
  .DOUT(bus_305dcfd3_), .DONE());
assign or_70dee808_u0=and_635d9962_u0|logicalMem_d0e13e1_we_delay0_u0;
assign and_635d9962_u0=bus_0aab59c9_&not_4794121a_u0;
endmodule



module resized_LH2_xy_stateVar_Out1PortEnable(bus_08bf0a8c_, bus_5fdb8633_, bus_0abc9c50_, bus_79cef798_, bus_52d26b67_);
input		bus_08bf0a8c_;
input		bus_5fdb8633_;
input		bus_0abc9c50_;
input		bus_79cef798_;
output		bus_52d26b67_;
reg		stateVar_Out1PortEnable_u4=1'h0;
assign bus_52d26b67_=stateVar_Out1PortEnable_u4;
always @(posedge bus_08bf0a8c_ or posedge bus_5fdb8633_)
begin
if (bus_5fdb8633_)
stateVar_Out1PortEnable_u4<=1'h0;
else if (bus_0abc9c50_)
stateVar_Out1PortEnable_u4<=bus_79cef798_;
end
endmodule



module resized_LH2_xy_simplememoryreferee_7c0f4a30_(bus_10a19532_, bus_5397d7e3_, bus_020ff5a4_, bus_06009997_, bus_7a5e2484_, bus_60ad4ce1_, bus_0309c2e0_, bus_0b593446_, bus_05ee34dd_, bus_56490b57_, bus_5b40276e_, bus_7aff8d40_, bus_19414a38_, bus_54364352_, bus_7a0b085e_, bus_180d93a2_, bus_05401935_, bus_736af7eb_, bus_04f85a99_, bus_50563d51_, bus_4687e307_, bus_307decb9_, bus_4686658d_, bus_13df4b68_);
input		bus_10a19532_;
input		bus_5397d7e3_;
input		bus_020ff5a4_;
input	[15:0]	bus_06009997_;
input		bus_7a5e2484_;
input	[15:0]	bus_60ad4ce1_;
input	[31:0]	bus_0309c2e0_;
input	[2:0]	bus_0b593446_;
input		bus_05ee34dd_;
input	[15:0]	bus_56490b57_;
input	[31:0]	bus_5b40276e_;
input	[2:0]	bus_7aff8d40_;
input		bus_19414a38_;
input	[31:0]	bus_54364352_;
input	[2:0]	bus_7a0b085e_;
output	[15:0]	bus_180d93a2_;
output	[31:0]	bus_05401935_;
output		bus_736af7eb_;
output		bus_04f85a99_;
output	[2:0]	bus_50563d51_;
output		bus_4687e307_;
output		bus_307decb9_;
output	[15:0]	bus_4686658d_;
output		bus_13df4b68_;
wire		and_56f1da31_u0;
reg		done_qual_u197_u0=1'h0;
wire		or_01217922_u0;
wire		or_2517a4f3_u0;
wire		not_1dc17be4_u0;
wire	[31:0]	mux_2b6f5aa7_u0;
wire		and_4186362e_u0;
wire	[15:0]	mux_1b60fd2a_u0;
reg		done_qual_u198_u0=1'h0;
wire		and_01ea51d8_u0;
wire		not_0e87bb35_u0;
wire		or_230435b1_u0;
reg		done_qual_u199_u0=1'h0;
wire		not_2fb6dd6d_u0;
wire		or_3db5ff28_u0;
wire		or_671226ad_u0;
assign and_56f1da31_u0=or_671226ad_u0&bus_020ff5a4_;
always @(posedge bus_10a19532_)
begin
if (bus_5397d7e3_)
done_qual_u197_u0<=1'h0;
else done_qual_u197_u0<=bus_19414a38_;
end
assign or_01217922_u0=bus_7a5e2484_|bus_05ee34dd_;
assign or_2517a4f3_u0=bus_19414a38_|done_qual_u197_u0;
assign bus_180d93a2_=mux_1b60fd2a_u0;
assign bus_05401935_=mux_2b6f5aa7_u0;
assign bus_736af7eb_=or_01217922_u0;
assign bus_04f85a99_=or_230435b1_u0;
assign bus_50563d51_=3'h1;
assign bus_4687e307_=and_56f1da31_u0;
assign bus_307decb9_=and_01ea51d8_u0;
assign bus_4686658d_=bus_06009997_;
assign bus_13df4b68_=and_4186362e_u0;
assign not_1dc17be4_u0=~bus_020ff5a4_;
assign mux_2b6f5aa7_u0=({32{bus_7a5e2484_}}&bus_0309c2e0_)|({32{bus_05ee34dd_}}&bus_5b40276e_)|({32{bus_19414a38_}}&bus_54364352_);
assign and_4186362e_u0=or_2517a4f3_u0&bus_020ff5a4_;
assign mux_1b60fd2a_u0=(bus_7a5e2484_)?bus_60ad4ce1_:bus_56490b57_;
always @(posedge bus_10a19532_)
begin
if (bus_5397d7e3_)
done_qual_u198_u0<=1'h0;
else done_qual_u198_u0<=bus_05ee34dd_;
end
assign and_01ea51d8_u0=or_3db5ff28_u0&bus_020ff5a4_;
assign not_0e87bb35_u0=~bus_020ff5a4_;
assign or_230435b1_u0=bus_7a5e2484_|bus_05ee34dd_|bus_19414a38_;
always @(posedge bus_10a19532_)
begin
if (bus_5397d7e3_)
done_qual_u199_u0<=1'h0;
else done_qual_u199_u0<=bus_7a5e2484_;
end
assign not_2fb6dd6d_u0=~bus_020ff5a4_;
assign or_3db5ff28_u0=bus_05ee34dd_|done_qual_u198_u0;
assign or_671226ad_u0=bus_7a5e2484_|done_qual_u199_u0;
endmodule


