// __  ___ __ ___  _ __   ___  ___ 
// \ \/ / '__/ _ \| '_ \ / _ \/ __|
//  >  <| | | (_) | | | | (_) \__ \
// /_/\_\_|  \___/|_| |_|\___/|___/
// 
// Xronos synthesizer version
// Run date: Thu 2 Nov 2017 13:58:31 +0000
// 

module image1_iunzip(Out2_DATA, Out1_RDY, Out2_RDY, Out1_ACK, Out1_COUNT, Out1_SEND, Out2_SEND, Out2_COUNT, CLK, RESET, In1_DATA, Out1_DATA, In1_COUNT, Out2_ACK, In1_ACK, In1_SEND);
output	[15:0]	Out2_DATA;
input		Out1_RDY;
input		Out2_RDY;
input		Out1_ACK;
output	[15:0]	Out1_COUNT;
wire		firstNPixels_go;
output		Out1_SEND;
output		Out2_SEND;
wire		firstNPixels_done;
wire		streamFun1_done;
wire		streamEndFun2_go;
output	[15:0]	Out2_COUNT;
wire		streamEndFun1_go;
wire		streamFun2_done;
input		CLK;
wire		streamEndFun2_done;
input		RESET;
input	[15:0]	In1_DATA;
output	[15:0]	Out1_DATA;
input	[15:0]	In1_COUNT;
input		Out2_ACK;
wire		streamEndFun1_done;
wire		streamFun2_go;
output		In1_ACK;
wire		streamFun1_go;
input		In1_SEND;
wire	[15:0]	bus_0b4f8702_;
wire		bus_6996ee9c_;
wire	[15:0]	bus_45f2eb26_;
wire		bus_09ba8778_;
wire	[1:0]	bus_713e8b32_;
wire	[31:0]	bus_412808a9_;
wire		bus_4b6527d6_;
wire	[2:0]	streamEndFun1_u3;
wire	[15:0]	streamEndFun1_u12;
wire	[31:0]	streamEndFun1_u5;
wire	[31:0]	streamEndFun1_u2;
wire		streamEndFun1_u4;
wire	[15:0]	streamEndFun1_u11;
wire		streamEndFun1;
wire		image1_iunzip_streamEndFun1_instance_DONE;
wire		streamEndFun1_u9;
wire		streamEndFun1_u0;
wire	[15:0]	streamEndFun1_u7;
wire		streamEndFun1_u10;
wire	[15:0]	streamEndFun1_u8;
wire	[2:0]	streamEndFun1_u6;
wire		streamEndFun1_u1;
wire	[1:0]	bus_0d633a7d_;
wire		bus_0eff1eb4_;
wire		or_7f062a31_u0;
wire		streamFun2;
wire	[15:0]	streamFun2_u13;
wire		streamFun2_u1;
wire	[31:0]	streamFun2_u2;
wire		streamFun2_u3;
wire	[31:0]	streamFun2_u4;
wire	[2:0]	streamFun2_u12;
wire		image1_iunzip_streamFun2_instance_DONE;
wire	[2:0]	streamFun2_u8;
wire	[31:0]	streamFun2_u10;
wire		streamFun2_u0;
wire		streamFun2_u14;
wire	[15:0]	streamFun2_u11;
wire		streamFun2_u15;
wire		streamFun2_u6;
wire		streamFun2_u9;
wire	[15:0]	streamFun2_u16;
wire	[31:0]	streamFun2_u7;
wire	[2:0]	streamFun2_u5;
wire		bus_79302887_;
wire		bus_028a7811_;
wire	[31:0]	bus_6bbd8c15_;
wire		or_7c8b174c_u0;
wire	[15:0]	or_403b04f2_u0;
wire	[31:0]	bus_6d8ec6c0_;
wire	[15:0]	bus_01bb560e_;
wire	[15:0]	bus_185cf169_;
wire	[2:0]	bus_3f0f2b61_;
wire	[15:0]	bus_1de509a3_;
wire		bus_2e00db39_;
wire		bus_438eba07_;
wire	[15:0]	bus_349fc2ad_;
wire		bus_380af87e_;
wire	[31:0]	bus_711ba866_;
wire		bus_3d439865_;
wire		bus_3c8caa47_;
wire	[15:0]	bus_5f260ad4_;
wire		bus_7818c025_;
wire		bus_0a070650_;
wire		streamFun1_u0;
wire	[2:0]	streamFun1_u5;
wire		streamFun1_u6;
wire		streamFun1_u1;
wire	[31:0]	streamFun1_u2;
wire		streamFun1_u3;
wire	[15:0]	streamFun1_u11;
wire		streamFun1_u14;
wire	[15:0]	streamFun1_u13;
wire	[31:0]	streamFun1_u10;
wire	[31:0]	streamFun1_u7;
wire		streamFun1_u16;
wire		streamFun1;
wire		streamFun1_u9;
wire	[2:0]	streamFun1_u12;
wire		image1_iunzip_streamFun1_instance_DONE;
wire	[31:0]	streamFun1_u4;
wire	[2:0]	streamFun1_u8;
wire	[15:0]	streamFun1_u15;
wire		or_77fce0a7_u0;
wire		bus_4d510363_;
wire	[31:0]	bus_59b1b34a_;
wire	[2:0]	bus_6aac9d02_;
wire	[15:0]	bus_56d7b0af_;
wire		bus_5b4fce35_;
wire		bus_4ef7394f_;
wire	[15:0]	bus_3f4ce93d_;
wire		bus_26adeb9f_;
wire	[15:0]	or_6a009060_u0;
wire	[15:0]	or_07ec3e80_u0;
wire		bus_0532da99_;
wire	[15:0]	or_26a54bd6_u0;
wire	[1:0]	scheduler_u86;
wire		scheduler;
wire		scheduler_u89;
wire		scheduler_u91;
wire	[2:0]	scheduler_u98;
wire	[31:0]	scheduler_u92;
wire		scheduler_u104;
wire		scheduler_u103;
wire		scheduler_u101;
wire		image1_iunzip_scheduler_instance_DONE;
wire	[1:0]	scheduler_u88;
wire		scheduler_u99;
wire		scheduler_u93;
wire		scheduler_u100;
wire		scheduler_u102;
wire		scheduler_u94;
wire	[15:0]	scheduler_u97;
wire		scheduler_u95;
wire		scheduler_u87;
wire	[31:0]	scheduler_u90;
wire	[31:0]	scheduler_u96;
wire	[31:0]	bus_592fb24a_;
wire		bus_4399e227_;
wire		bus_68afb47e_;
wire	[15:0]	bus_73bd858d_;
wire		bus_1604219b_;
wire	[2:0]	bus_7a726660_;
wire	[15:0]	bus_4ba2e658_;
wire		bus_394326ad_;
wire		bus_5857bbf3_;
wire		bus_6204046f_;
wire	[15:0]	bus_0c649092_;
wire	[15:0]	bus_6d3e7bde_;
wire		bus_4cc7a537_;
wire	[15:0]	streamEndFun2_u8;
wire	[31:0]	streamEndFun2_u5;
wire		streamEndFun2_u0;
wire		streamEndFun2_u1;
wire	[15:0]	streamEndFun2_u7;
wire	[15:0]	streamEndFun2_u11;
wire	[2:0]	streamEndFun2_u3;
wire	[31:0]	streamEndFun2_u2;
wire		streamEndFun2;
wire	[15:0]	streamEndFun2_u12;
wire	[2:0]	streamEndFun2_u6;
wire		streamEndFun2_u9;
wire		streamEndFun2_u4;
wire		streamEndFun2_u10;
wire		image1_iunzip_streamEndFun2_instance_DONE;
wire		bus_71ee2f20_;
wire	[15:0]	firstNPixels_u6;
wire		firstNPixels_u8;
wire	[2:0]	firstNPixels_u3;
wire		firstNPixels_u4;
wire		firstNPixels_u1;
wire		image1_iunzip_firstNPixels_instance_DONE;
wire	[2:0]	firstNPixels_u7;
wire		firstNPixels;
wire	[31:0]	firstNPixels_u2;
wire	[31:0]	firstNPixels_u9;
wire	[2:0]	firstNPixels_u10;
wire	[31:0]	firstNPixels_u0;
wire	[31:0]	firstNPixels_u5;
wire		bus_1066ab06_;
wire		bus_225c3717_;
wire	[15:0]	bus_32560469_;
wire		bus_6b5b6b3c_;
wire	[15:0]	bus_0cf04c6c_;
wire	[15:0]	bus_3c871d5b_;
wire		bus_05e31049_;
wire	[15:0]	bus_52b719e4_;
wire		bus_3b62cf1f_;
wire	[2:0]	bus_4b0b58ac_;
wire		bus_1e395c9f_;
wire	[15:0]	bus_628ee2f9_;
wire	[31:0]	bus_0d379228_;
wire		bus_08315480_;
assign Out2_DATA=or_403b04f2_u0;
assign Out1_COUNT=or_26a54bd6_u0;
assign firstNPixels_go=scheduler_u99;
assign Out1_SEND=or_77fce0a7_u0;
assign Out2_SEND=or_7c8b174c_u0;
assign firstNPixels_done=bus_0eff1eb4_;
assign streamFun1_done=bus_028a7811_;
assign streamEndFun2_go=scheduler_u102;
assign Out2_COUNT=or_6a009060_u0;
assign streamEndFun1_go=scheduler_u104;
assign streamFun2_done=bus_4b6527d6_;
assign streamEndFun2_done=bus_26adeb9f_;
assign Out1_DATA=or_07ec3e80_u0;
assign streamEndFun1_done=bus_0a070650_;
assign streamFun2_go=scheduler_u101;
assign In1_ACK=or_7f062a31_u0;
assign streamFun1_go=scheduler_u100;
image1_iunzip_structuralmemory_590a638a_ image1_iunzip_structuralmemory_590a638a__1(.CLK_u2(CLK), 
  .bus_1e163efd_(bus_5857bbf3_), .bus_4e2d7f14_(32'h1), .bus_582a5b58_(3'h1), .bus_74db3565_(bus_4d510363_), 
  .bus_593523a5_(bus_592fb24a_), .bus_32f6c133_(3'h1), .bus_5f8c7c67_(bus_1604219b_), 
  .bus_70d2a891_(bus_68afb47e_), .bus_2906b104_(bus_73bd858d_), .bus_0b4f8702_(bus_0b4f8702_), 
  .bus_09ba8778_(bus_09ba8778_), .bus_45f2eb26_(bus_45f2eb26_), .bus_6996ee9c_(bus_6996ee9c_));
image1_iunzip_stateVar_fsmOldState_image1_iunzip image1_iunzip_stateVar_fsmOldState_image1_iunzip_1(.bus_1d4c8b6d_(CLK), 
  .bus_06f0cc30_(bus_5857bbf3_), .bus_1ca24d20_(scheduler), .bus_65dd6bff_(scheduler_u86), 
  .bus_713e8b32_(bus_713e8b32_));
image1_iunzip_stateVar_consumed image1_iunzip_stateVar_consumed_1(.bus_7118581b_(CLK), 
  .bus_146858d2_(bus_5857bbf3_), .bus_5ccce527_(firstNPixels), .bus_395fdddb_(firstNPixels_u0), 
  .bus_382b6c3a_(streamFun1_u1), .bus_2d19da07_(streamFun1_u2), .bus_67c9cda4_(streamFun2_u1), 
  .bus_150154ba_(streamFun2_u2), .bus_412808a9_(bus_412808a9_));
assign bus_4b6527d6_=image1_iunzip_streamFun2_instance_DONE&{1{image1_iunzip_streamFun2_instance_DONE}};
image1_iunzip_streamEndFun1 image1_iunzip_streamEndFun1_instance(.CLK(CLK), .RESET(bus_5857bbf3_), 
  .GO(streamEndFun1_go), .port_3927e736_(bus_79302887_), .port_1f3f2d39_(bus_1066ab06_), 
  .port_1df607d4_(bus_32560469_), .port_7b58ab67_(bus_7818c025_), .port_129b8bb2_(bus_349fc2ad_), 
  .DONE(image1_iunzip_streamEndFun1_instance_DONE), .RESULT(streamEndFun1), .RESULT_u740(streamEndFun1_u0), 
  .RESULT_u741(streamEndFun1_u1), .RESULT_u742(streamEndFun1_u2), .RESULT_u743(streamEndFun1_u3), 
  .RESULT_u744(streamEndFun1_u4), .RESULT_u745(streamEndFun1_u5), .RESULT_u746(streamEndFun1_u6), 
  .RESULT_u747(streamEndFun1_u7), .RESULT_u748(streamEndFun1_u8), .RESULT_u749(streamEndFun1_u9), 
  .RESULT_u750(streamEndFun1_u10), .RESULT_u751(streamEndFun1_u11), .RESULT_u752(streamEndFun1_u12));
image1_iunzip_stateVar_fsmState_image1_iunzip image1_iunzip_stateVar_fsmState_image1_iunzip_1(.bus_4c915309_(CLK), 
  .bus_2d7bb642_(bus_5857bbf3_), .bus_02e4d33b_(scheduler_u87), .bus_3412b614_(scheduler_u88), 
  .bus_0d633a7d_(bus_0d633a7d_));
assign bus_0eff1eb4_=image1_iunzip_firstNPixels_instance_DONE&{1{image1_iunzip_firstNPixels_instance_DONE}};
assign or_7f062a31_u0=streamFun1_u16|streamFun2_u15|scheduler_u103;
image1_iunzip_streamFun2 image1_iunzip_streamFun2_instance(.CLK(CLK), .RESET(bus_5857bbf3_), 
  .GO(streamFun2_go), .port_4da7fcea_(bus_79302887_), .port_5ec353a6_(bus_412808a9_), 
  .port_001ed422_(bus_3c8caa47_), .port_08ebfbc1_(bus_01bb560e_), .port_45273060_(bus_05e31049_), 
  .port_221c496a_(bus_0cf04c6c_), .port_0ebd1361_(bus_05e31049_), .port_587fd1a5_(In1_DATA), 
  .DONE(image1_iunzip_streamFun2_instance_DONE), .RESULT(streamFun2), .RESULT_u753(streamFun2_u0), 
  .RESULT_u754(streamFun2_u1), .RESULT_u755(streamFun2_u2), .RESULT_u763(streamFun2_u3), 
  .RESULT_u764(streamFun2_u4), .RESULT_u765(streamFun2_u5), .RESULT_u756(streamFun2_u6), 
  .RESULT_u757(streamFun2_u7), .RESULT_u758(streamFun2_u8), .RESULT_u759(streamFun2_u9), 
  .RESULT_u760(streamFun2_u10), .RESULT_u761(streamFun2_u11), .RESULT_u762(streamFun2_u12), 
  .RESULT_u766(streamFun2_u13), .RESULT_u767(streamFun2_u14), .RESULT_u768(streamFun2_u15), 
  .RESULT_u769(streamFun2_u16));
image1_iunzip_stateVar_midPoint image1_iunzip_stateVar_midPoint_1(.bus_676a86b4_(CLK), 
  .bus_7f9b1e16_(bus_5857bbf3_), .bus_6d113f7e_(streamFun1), .bus_79b19529_(1'h0), 
  .bus_196aa05d_(streamFun2), .bus_5894ff4e_(1'h0), .bus_4ddfe8ac_(streamEndFun1), 
  .bus_56ab03e3_(1'h0), .bus_3b63cd45_(streamEndFun2), .bus_4ba5b0a8_(1'h0), .bus_79302887_(bus_79302887_));
assign bus_028a7811_=image1_iunzip_streamFun1_instance_DONE&{1{image1_iunzip_streamFun1_instance_DONE}};
image1_iunzip_stateVar_In1TokenIndex image1_iunzip_stateVar_In1TokenIndex_1(.bus_00a6f1a7_(CLK), 
  .bus_05ce656d_(bus_5857bbf3_), .bus_69335eb2_(scheduler_u89), .bus_28bc525f_(scheduler_u90), 
  .bus_6bbd8c15_(bus_6bbd8c15_));
assign or_7c8b174c_u0=streamFun2_u14|streamEndFun1_u10|streamEndFun2_u10;
assign or_403b04f2_u0=streamFun2_u13|streamEndFun1_u8|streamEndFun2_u8;
image1_iunzip_stateVar_In1MaxTokenIndex image1_iunzip_stateVar_In1MaxTokenIndex_1(.bus_022df17c_(CLK), 
  .bus_1facd4e4_(bus_5857bbf3_), .bus_4a9eda6d_(scheduler_u91), .bus_5e278fb9_({scheduler_u92[31:2], 1'b0, scheduler_u92[0]}), 
  .bus_6d8ec6c0_(bus_6d8ec6c0_));
image1_iunzip_simplememoryreferee_0b0f52d7_ image1_iunzip_simplememoryreferee_0b0f52d7__1(.bus_29cdd1f8_(CLK), 
  .bus_6b72c155_(bus_5857bbf3_), .bus_3c855b7b_(bus_4cc7a537_), .bus_20f0729f_(bus_0c649092_), 
  .bus_5b77758f_(streamFun1_u3), .bus_5b45fa2c_(streamFun1_u4), .bus_0964b8c9_(3'h1), 
  .bus_37539c61_(streamFun2_u3), .bus_1daba9ee_(streamFun2_u4), .bus_0e50a633_(3'h1), 
  .bus_6d9883cb_(streamEndFun1_u4), .bus_5525d2cf_(streamEndFun1_u5), .bus_5038a20c_(3'h1), 
  .bus_267b146b_(streamEndFun2_u4), .bus_67995a05_(streamEndFun2_u5), .bus_5fbad179_(3'h1), 
  .bus_5f260ad4_(bus_5f260ad4_), .bus_711ba866_(bus_711ba866_), .bus_3d439865_(bus_3d439865_), 
  .bus_2e00db39_(bus_2e00db39_), .bus_3f0f2b61_(bus_3f0f2b61_), .bus_1de509a3_(bus_1de509a3_), 
  .bus_438eba07_(bus_438eba07_), .bus_01bb560e_(bus_01bb560e_), .bus_3c8caa47_(bus_3c8caa47_), 
  .bus_349fc2ad_(bus_349fc2ad_), .bus_7818c025_(bus_7818c025_), .bus_185cf169_(bus_185cf169_), 
  .bus_380af87e_(bus_380af87e_));
assign bus_0a070650_=image1_iunzip_streamEndFun1_instance_DONE&{1{image1_iunzip_streamEndFun1_instance_DONE}};
image1_iunzip_streamFun1 image1_iunzip_streamFun1_instance(.CLK(CLK), .RESET(bus_5857bbf3_), 
  .GO(streamFun1_go), .port_4691c47d_(bus_79302887_), .port_0289ded9_(bus_412808a9_), 
  .port_7ab2bf13_(bus_438eba07_), .port_6ecc5cde_(bus_1de509a3_), .port_635f8008_(bus_225c3717_), 
  .port_747b457f_(bus_3c871d5b_), .port_1d854cce_(bus_225c3717_), .port_01e6d96a_(In1_DATA), 
  .DONE(image1_iunzip_streamFun1_instance_DONE), .RESULT(streamFun1), .RESULT_u770(streamFun1_u0), 
  .RESULT_u771(streamFun1_u1), .RESULT_u772(streamFun1_u2), .RESULT_u780(streamFun1_u3), 
  .RESULT_u781(streamFun1_u4), .RESULT_u782(streamFun1_u5), .RESULT_u773(streamFun1_u6), 
  .RESULT_u774(streamFun1_u7), .RESULT_u775(streamFun1_u8), .RESULT_u776(streamFun1_u9), 
  .RESULT_u777(streamFun1_u10), .RESULT_u778(streamFun1_u11), .RESULT_u779(streamFun1_u12), 
  .RESULT_u783(streamFun1_u13), .RESULT_u784(streamFun1_u14), .RESULT_u785(streamFun1_u15), 
  .RESULT_u786(streamFun1_u16));
assign or_77fce0a7_u0=streamFun1_u14|streamEndFun1_u9|streamEndFun2_u9;
image1_iunzip_simplememoryreferee_4f4a8814_ image1_iunzip_simplememoryreferee_4f4a8814__1(.bus_6a794fd6_(CLK), 
  .bus_561f7191_(bus_5857bbf3_), .bus_495872da_(bus_09ba8778_), .bus_220964f4_(bus_0b4f8702_), 
  .bus_31862682_(firstNPixels_u8), .bus_0040cf15_(32'h1), .bus_5ccabeca_(3'h1), 
  .bus_56d7b0af_(bus_56d7b0af_), .bus_59b1b34a_(bus_59b1b34a_), .bus_5b4fce35_(bus_5b4fce35_), 
  .bus_4d510363_(bus_4d510363_), .bus_6aac9d02_(bus_6aac9d02_), .bus_3f4ce93d_(bus_3f4ce93d_), 
  .bus_4ef7394f_(bus_4ef7394f_));
assign bus_26adeb9f_=image1_iunzip_streamEndFun2_instance_DONE&{1{image1_iunzip_streamEndFun2_instance_DONE}};
assign or_6a009060_u0=streamFun2_u16|streamEndFun1_u12|streamEndFun2_u12;
assign or_07ec3e80_u0=streamFun1_u15|streamEndFun1_u11|streamEndFun2_u11;
image1_iunzip_Kicker_22 image1_iunzip_Kicker_22_1(.CLK(CLK), .RESET(bus_5857bbf3_), 
  .bus_0532da99_(bus_0532da99_));
assign or_26a54bd6_u0=streamFun1_u13|streamEndFun1_u7|streamEndFun2_u7;
image1_iunzip_scheduler image1_iunzip_scheduler_instance(.CLK(CLK), .RESET(bus_5857bbf3_), 
  .GO(bus_0532da99_), .port_18e00d02_(bus_713e8b32_), .port_7b9868d2_(bus_0d633a7d_), 
  .port_5b5cde36_(bus_6bbd8c15_), .port_7a3e2d5e_(bus_6d8ec6c0_), .port_2b235147_(bus_412808a9_), 
  .port_30bf0bb1_(bus_4399e227_), .port_2d451d49_(Out1_RDY), .port_01ffd1e5_(Out2_RDY), 
  .port_6c59504e_(streamEndFun1_done), .port_7dc7ca1e_(In1_DATA), .port_2f06a0cc_(streamFun1_done), 
  .port_2cc0cc2a_(In1_SEND), .port_65a60be6_(firstNPixels_done), .port_0312d0b7_(streamEndFun2_done), 
  .port_4fbbb17b_(streamFun2_done), .DONE(image1_iunzip_scheduler_instance_DONE), 
  .RESULT(scheduler), .RESULT_u787(scheduler_u86), .RESULT_u788(scheduler_u87), 
  .RESULT_u789(scheduler_u88), .RESULT_u790(scheduler_u89), .RESULT_u791(scheduler_u90), 
  .RESULT_u792(scheduler_u91), .RESULT_u793(scheduler_u92), .RESULT_u794(scheduler_u93), 
  .RESULT_u795(scheduler_u94), .RESULT_u796(scheduler_u95), .RESULT_u797(scheduler_u96), 
  .RESULT_u798(scheduler_u97), .RESULT_u799(scheduler_u98), .RESULT_u800(scheduler_u99), 
  .RESULT_u801(scheduler_u100), .RESULT_u802(scheduler_u101), .RESULT_u803(scheduler_u102), 
  .RESULT_u804(scheduler_u103), .RESULT_u805(scheduler_u104));
image1_iunzip_simplememoryreferee_3f8b2b7e_ image1_iunzip_simplememoryreferee_3f8b2b7e__1(.bus_4fdc6d9e_(CLK), 
  .bus_16db627b_(bus_5857bbf3_), .bus_5c6b1ef6_(bus_6996ee9c_), .bus_7e5a1f5a_(bus_45f2eb26_), 
  .bus_220ac51f_(firstNPixels_u1), .bus_77abea3c_(32'h0), .bus_55f9978e_(3'h1), 
  .bus_192ef9bb_(scheduler_u95), .bus_26fb90a8_(scheduler_u97), .bus_5ac8d702_(scheduler_u96), 
  .bus_5fd8a7cf_(3'h1), .bus_73bd858d_(bus_73bd858d_), .bus_592fb24a_(bus_592fb24a_), 
  .bus_68afb47e_(bus_68afb47e_), .bus_1604219b_(bus_1604219b_), .bus_7a726660_(bus_7a726660_), 
  .bus_4ba2e658_(bus_4ba2e658_), .bus_394326ad_(bus_394326ad_), .bus_4399e227_(bus_4399e227_));
image1_iunzip_globalreset_physical_0787df71_ image1_iunzip_globalreset_physical_0787df71__1(.bus_137e2708_(CLK), 
  .bus_19659027_(RESET), .bus_5857bbf3_(bus_5857bbf3_));
image1_iunzip_structuralmemory_224e8538_ image1_iunzip_structuralmemory_224e8538__1(.CLK_u3(CLK), 
  .bus_44b4fa91_(bus_5857bbf3_), .bus_0f1d20b4_(bus_0d379228_), .bus_625040d8_(3'h1), 
  .bus_38cab4e5_(bus_3b62cf1f_), .bus_1f7bdd2e_(bus_1e395c9f_), .bus_4944043d_(bus_628ee2f9_), 
  .bus_2448127a_(bus_711ba866_), .bus_016e260c_(3'h1), .bus_25f12fe5_(bus_2e00db39_), 
  .bus_6d3e7bde_(bus_6d3e7bde_), .bus_6204046f_(bus_6204046f_), .bus_0c649092_(bus_0c649092_), 
  .bus_4cc7a537_(bus_4cc7a537_));
image1_iunzip_streamEndFun2 image1_iunzip_streamEndFun2_instance(.CLK(CLK), .RESET(bus_5857bbf3_), 
  .GO(streamEndFun2_go), .port_63ac392a_(bus_79302887_), .port_4739a893_(bus_08315480_), 
  .port_2068be2c_(bus_52b719e4_), .port_1e8c51ba_(bus_380af87e_), .port_177ce6b0_(bus_185cf169_), 
  .DONE(image1_iunzip_streamEndFun2_instance_DONE), .RESULT(streamEndFun2), .RESULT_u806(streamEndFun2_u0), 
  .RESULT_u807(streamEndFun2_u1), .RESULT_u808(streamEndFun2_u2), .RESULT_u809(streamEndFun2_u3), 
  .RESULT_u810(streamEndFun2_u4), .RESULT_u811(streamEndFun2_u5), .RESULT_u812(streamEndFun2_u6), 
  .RESULT_u813(streamEndFun2_u7), .RESULT_u814(streamEndFun2_u8), .RESULT_u815(streamEndFun2_u9), 
  .RESULT_u816(streamEndFun2_u10), .RESULT_u817(streamEndFun2_u11), .RESULT_u818(streamEndFun2_u12));
image1_iunzip_stateVar_In1PortEnable image1_iunzip_stateVar_In1PortEnable_1(.bus_6b4f1791_(CLK), 
  .bus_7b3d8b32_(bus_5857bbf3_), .bus_1712d9e1_(scheduler_u93), .bus_1301d8aa_(scheduler_u94), 
  .bus_71ee2f20_(bus_71ee2f20_));
image1_iunzip_firstNPixels image1_iunzip_firstNPixels_instance(.CLK(CLK), .RESET(bus_5857bbf3_), 
  .GO(firstNPixels_go), .port_0e7ec45d_(bus_412808a9_), .port_30f2a2a5_(bus_394326ad_), 
  .port_58472f4a_(bus_4ba2e658_), .port_10601e70_(bus_6b5b6b3c_), .port_328b25f5_(bus_4ef7394f_), 
  .port_33fbecb1_(bus_3f4ce93d_), .DONE(image1_iunzip_firstNPixels_instance_DONE), 
  .RESULT(firstNPixels), .RESULT_u819(firstNPixels_u0), .RESULT_u827(firstNPixels_u1), 
  .RESULT_u828(firstNPixels_u2), .RESULT_u829(firstNPixels_u3), .RESULT_u820(firstNPixels_u4), 
  .RESULT_u821(firstNPixels_u5), .RESULT_u822(firstNPixels_u6), .RESULT_u823(firstNPixels_u7), 
  .RESULT_u824(firstNPixels_u8), .RESULT_u825(firstNPixels_u9), .RESULT_u826(firstNPixels_u10));
image1_iunzip_simplememoryreferee_12559ca8_ image1_iunzip_simplememoryreferee_12559ca8__1(.bus_34d6401e_(CLK), 
  .bus_2c677a40_(bus_5857bbf3_), .bus_61602789_(bus_6204046f_), .bus_520a81dd_(bus_6d3e7bde_), 
  .bus_4f242077_(firstNPixels_u4), .bus_56e7637f_(firstNPixels_u6), .bus_2414a2f1_({31'b0, firstNPixels_u5[0]}), 
  .bus_4906a1e5_(3'h1), .bus_0cb5957a_(streamFun1_u6), .bus_4c5426bf_(streamFun1_u9), 
  .bus_4034cf94_(streamFun1_u11), .bus_12ed058a_(streamFun1_u10), .bus_50e7e991_(3'h1), 
  .bus_4f572e1e_(streamFun2_u6), .bus_20b4c307_(streamFun2_u9), .bus_32b5a413_(streamFun2_u11), 
  .bus_4b85717f_(streamFun2_u10), .bus_3181df50_(3'h1), .bus_2f2a289d_(streamEndFun1_u1), 
  .bus_25006614_(streamEndFun1_u2), .bus_4d322080_(3'h1), .bus_77aca28c_(streamEndFun2_u1), 
  .bus_6af53624_(streamEndFun2_u2), .bus_0a775a74_(3'h1), .bus_628ee2f9_(bus_628ee2f9_), 
  .bus_0d379228_(bus_0d379228_), .bus_1e395c9f_(bus_1e395c9f_), .bus_3b62cf1f_(bus_3b62cf1f_), 
  .bus_4b0b58ac_(bus_4b0b58ac_), .bus_6b5b6b3c_(bus_6b5b6b3c_), .bus_3c871d5b_(bus_3c871d5b_), 
  .bus_225c3717_(bus_225c3717_), .bus_0cf04c6c_(bus_0cf04c6c_), .bus_05e31049_(bus_05e31049_), 
  .bus_32560469_(bus_32560469_), .bus_1066ab06_(bus_1066ab06_), .bus_52b719e4_(bus_52b719e4_), 
  .bus_08315480_(bus_08315480_));
endmodule



module image1_iunzip_forge_memory_2x16_6(CLK, ENA, WEA, DINA, ENB, ADDRA, ADDRB, DOUTA, DOUTB, DONEA, DONEB);
input		CLK;
input		ENA;
input		WEA;
input	[15:0]	DINA;
input		ENB;
input	[31:0]	ADDRA;
input	[31:0]	ADDRB;
output	[15:0]	DOUTA;
output	[15:0]	DOUTB;
output		DONEA;
output		DONEB;
wire		wea_0;
wire	[15:0]	pre_douta_0;
wire	[15:0]	pre_doutb_0;
reg		wea_done;
reg		rea_done;
reg	[15:0]	mux_outa;
reg	[15:0]	mux_outb;
assign wea_0=WEA;
always @(posedge CLK)
begin
wea_done<=WEA;
end
assign DONEA=rea_done|wea_done;
always @(posedge CLK)
begin
end
assign DONEB=ENB;
always @(pre_douta_0)
begin
mux_outa<=pre_douta_0;
end
assign DOUTA=mux_outa;
always @(pre_doutb_0)
begin
mux_outb<=pre_doutb_0;
end
assign DOUTB=mux_outb;
// Memory array element: COL: 0, ROW: 0
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_0(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[0]), .SPO(pre_douta_0[0]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[0]));
// Memory array element: COL: 0, ROW: 1
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_1(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[1]), .SPO(pre_douta_0[1]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[1]));
// Memory array element: COL: 0, ROW: 2
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_2(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[2]), .SPO(pre_douta_0[2]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[2]));
// Memory array element: COL: 0, ROW: 3
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_3(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[3]), .SPO(pre_douta_0[3]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[3]));
// Memory array element: COL: 0, ROW: 4
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_4(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[4]), .SPO(pre_douta_0[4]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[4]));
// Memory array element: COL: 0, ROW: 5
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_5(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[5]), .SPO(pre_douta_0[5]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[5]));
// Memory array element: COL: 0, ROW: 6
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_6(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[6]), .SPO(pre_douta_0[6]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[6]));
// Memory array element: COL: 0, ROW: 7
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_7(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[7]), .SPO(pre_douta_0[7]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[7]));
// Memory array element: COL: 0, ROW: 8
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_8(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[8]), .SPO(pre_douta_0[8]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[8]));
// Memory array element: COL: 0, ROW: 9
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_9(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[9]), .SPO(pre_douta_0[9]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[9]));
// Memory array element: COL: 0, ROW: 10
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_10(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[10]), .SPO(pre_douta_0[10]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[10]));
// Memory array element: COL: 0, ROW: 11
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_11(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[11]), .SPO(pre_douta_0[11]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[11]));
// Memory array element: COL: 0, ROW: 12
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_12(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[12]), .SPO(pre_douta_0[12]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[12]));
// Memory array element: COL: 0, ROW: 13
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_13(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[13]), .SPO(pre_douta_0[13]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[13]));
// Memory array element: COL: 0, ROW: 14
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_14(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[14]), .SPO(pre_douta_0[14]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[14]));
// Memory array element: COL: 0, ROW: 15
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_15(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[15]), .SPO(pre_douta_0[15]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[15]));
endmodule



module image1_iunzip_structuralmemory_590a638a_(CLK_u2, bus_1e163efd_, bus_4e2d7f14_, bus_582a5b58_, bus_74db3565_, bus_593523a5_, bus_32f6c133_, bus_5f8c7c67_, bus_70d2a891_, bus_2906b104_, bus_0b4f8702_, bus_09ba8778_, bus_45f2eb26_, bus_6996ee9c_);
input		CLK_u2;
input		bus_1e163efd_;
input	[31:0]	bus_4e2d7f14_;
input	[2:0]	bus_582a5b58_;
input		bus_74db3565_;
input	[31:0]	bus_593523a5_;
input	[2:0]	bus_32f6c133_;
input		bus_5f8c7c67_;
input		bus_70d2a891_;
input	[15:0]	bus_2906b104_;
output	[15:0]	bus_0b4f8702_;
output		bus_09ba8778_;
output	[15:0]	bus_45f2eb26_;
output		bus_6996ee9c_;
reg		logicalMem_a2e6c14_we_delay0_u0=1'h0;
wire		and_17700a68_u0;
wire		not_12c4497f_u0;
wire	[15:0]	bus_46a4089f_;
wire	[15:0]	bus_424a2dda_;
wire		or_55b98be7_u0;
wire		or_7c197906_u0;
assign bus_0b4f8702_=bus_46a4089f_;
assign bus_09ba8778_=bus_74db3565_;
assign bus_45f2eb26_=bus_424a2dda_;
assign bus_6996ee9c_=or_55b98be7_u0;
always @(posedge CLK_u2 or posedge bus_1e163efd_)
begin
if (bus_1e163efd_)
logicalMem_a2e6c14_we_delay0_u0<=1'h0;
else logicalMem_a2e6c14_we_delay0_u0<=bus_70d2a891_;
end
assign and_17700a68_u0=bus_5f8c7c67_&not_12c4497f_u0;
assign not_12c4497f_u0=~bus_70d2a891_;
image1_iunzip_forge_memory_2x16_6 image1_iunzip_forge_memory_2x16_6_instance0(.CLK(CLK_u2), 
  .ENA(or_7c197906_u0), .WEA(bus_70d2a891_), .DINA(bus_2906b104_), .ADDRA(bus_593523a5_), 
  .DOUTA(bus_424a2dda_), .DONEA(), .ENB(bus_74db3565_), .ADDRB(32'h1), .DOUTB(bus_46a4089f_), 
  .DONEB());
assign or_55b98be7_u0=and_17700a68_u0|logicalMem_a2e6c14_we_delay0_u0;
assign or_7c197906_u0=bus_5f8c7c67_|bus_70d2a891_;
endmodule



module image1_iunzip_endianswapper_55945173_(endianswapper_55945173_in, endianswapper_55945173_out);
input	[1:0]	endianswapper_55945173_in;
output	[1:0]	endianswapper_55945173_out;
assign endianswapper_55945173_out=endianswapper_55945173_in;
endmodule



module image1_iunzip_endianswapper_12ad75e2_(endianswapper_12ad75e2_in, endianswapper_12ad75e2_out);
input	[1:0]	endianswapper_12ad75e2_in;
output	[1:0]	endianswapper_12ad75e2_out;
assign endianswapper_12ad75e2_out=endianswapper_12ad75e2_in;
endmodule



module image1_iunzip_stateVar_fsmOldState_image1_iunzip(bus_1d4c8b6d_, bus_06f0cc30_, bus_1ca24d20_, bus_65dd6bff_, bus_713e8b32_);
input		bus_1d4c8b6d_;
input		bus_06f0cc30_;
input		bus_1ca24d20_;
input	[1:0]	bus_65dd6bff_;
output	[1:0]	bus_713e8b32_;
wire	[1:0]	endianswapper_55945173_out;
reg	[1:0]	stateVar_fsmOldState_image1_iunzip_u0=2'h0;
wire	[1:0]	endianswapper_12ad75e2_out;
image1_iunzip_endianswapper_55945173_ image1_iunzip_endianswapper_55945173__1(.endianswapper_55945173_in(bus_65dd6bff_), 
  .endianswapper_55945173_out(endianswapper_55945173_out));
always @(posedge bus_1d4c8b6d_ or posedge bus_06f0cc30_)
begin
if (bus_06f0cc30_)
stateVar_fsmOldState_image1_iunzip_u0<=2'h0;
else if (bus_1ca24d20_)
stateVar_fsmOldState_image1_iunzip_u0<=endianswapper_55945173_out;
end
assign bus_713e8b32_=endianswapper_12ad75e2_out;
image1_iunzip_endianswapper_12ad75e2_ image1_iunzip_endianswapper_12ad75e2__1(.endianswapper_12ad75e2_in(stateVar_fsmOldState_image1_iunzip_u0), 
  .endianswapper_12ad75e2_out(endianswapper_12ad75e2_out));
endmodule



module image1_iunzip_endianswapper_5e8c9437_(endianswapper_5e8c9437_in, endianswapper_5e8c9437_out);
input	[31:0]	endianswapper_5e8c9437_in;
output	[31:0]	endianswapper_5e8c9437_out;
assign endianswapper_5e8c9437_out=endianswapper_5e8c9437_in;
endmodule



module image1_iunzip_endianswapper_10599ef5_(endianswapper_10599ef5_in, endianswapper_10599ef5_out);
input	[31:0]	endianswapper_10599ef5_in;
output	[31:0]	endianswapper_10599ef5_out;
assign endianswapper_10599ef5_out=endianswapper_10599ef5_in;
endmodule



module image1_iunzip_stateVar_consumed(bus_7118581b_, bus_146858d2_, bus_5ccce527_, bus_395fdddb_, bus_382b6c3a_, bus_2d19da07_, bus_67c9cda4_, bus_150154ba_, bus_412808a9_);
input		bus_7118581b_;
input		bus_146858d2_;
input		bus_5ccce527_;
input	[31:0]	bus_395fdddb_;
input		bus_382b6c3a_;
input	[31:0]	bus_2d19da07_;
input		bus_67c9cda4_;
input	[31:0]	bus_150154ba_;
output	[31:0]	bus_412808a9_;
reg	[31:0]	stateVar_consumed_u2=32'h0;
wire	[31:0]	mux_35538a7b_u0;
wire	[31:0]	endianswapper_5e8c9437_out;
wire	[31:0]	endianswapper_10599ef5_out;
wire		or_4956ddf8_u0;
always @(posedge bus_7118581b_ or posedge bus_146858d2_)
begin
if (bus_146858d2_)
stateVar_consumed_u2<=32'h0;
else if (or_4956ddf8_u0)
stateVar_consumed_u2<=endianswapper_5e8c9437_out;
end
assign mux_35538a7b_u0=({32{bus_5ccce527_}}&bus_395fdddb_)|({32{bus_382b6c3a_}}&bus_2d19da07_)|({32{bus_67c9cda4_}}&bus_150154ba_);
assign bus_412808a9_=endianswapper_10599ef5_out;
image1_iunzip_endianswapper_5e8c9437_ image1_iunzip_endianswapper_5e8c9437__1(.endianswapper_5e8c9437_in(mux_35538a7b_u0), 
  .endianswapper_5e8c9437_out(endianswapper_5e8c9437_out));
image1_iunzip_endianswapper_10599ef5_ image1_iunzip_endianswapper_10599ef5__1(.endianswapper_10599ef5_in(stateVar_consumed_u2), 
  .endianswapper_10599ef5_out(endianswapper_10599ef5_out));
assign or_4956ddf8_u0=bus_5ccce527_|bus_382b6c3a_|bus_67c9cda4_;
endmodule



module image1_iunzip_streamEndFun1(CLK, RESET, GO, port_3927e736_, port_1f3f2d39_, port_1df607d4_, port_7b58ab67_, port_129b8bb2_, RESULT, RESULT_u740, RESULT_u741, RESULT_u742, RESULT_u743, RESULT_u744, RESULT_u745, RESULT_u746, RESULT_u747, RESULT_u748, RESULT_u749, RESULT_u750, RESULT_u751, RESULT_u752, DONE);
input		CLK;
input		RESET;
input		GO;
input		port_3927e736_;
input		port_1f3f2d39_;
input	[15:0]	port_1df607d4_;
input		port_7b58ab67_;
input	[15:0]	port_129b8bb2_;
output		RESULT;
output		RESULT_u740;
output		RESULT_u741;
output	[31:0]	RESULT_u742;
output	[2:0]	RESULT_u743;
output		RESULT_u744;
output	[31:0]	RESULT_u745;
output	[2:0]	RESULT_u746;
output	[15:0]	RESULT_u747;
output	[15:0]	RESULT_u748;
output		RESULT_u749;
output		RESULT_u750;
output	[15:0]	RESULT_u751;
output	[15:0]	RESULT_u752;
output		DONE;
wire	[31:0]	add;
wire		and_u1310_u0;
wire	[8:0]	subtract;
wire		greaterThanEqualTo;
wire signed	[8:0]	greaterThanEqualTo_a_signed;
wire signed	[8:0]	greaterThanEqualTo_b_signed;
wire		not_u252_u0;
wire		and_u1311_u0;
wire		and_u1312_u0;
wire	[8:0]	subtract_u0;
wire		and_u1313_u0;
wire		and_u1314_u0;
wire	[8:0]	mux_u80;
wire	[31:0]	add_u24;
wire		and_u1315_u0;
wire		and_u1317_u0;
wire	[16:0]	add_u25;
wire	[15:0]	subtract_u1;
wire	[15:0]	simplePinWrite;
wire	[15:0]	simplePinWrite_u212;
wire		simplePinWrite_u213;
wire	[15:0]	simplePinWrite_u214;
wire		simplePinWrite_u215;
wire	[15:0]	simplePinWrite_u216;
wire	[31:0]	mux_u81_u0;
wire		or_u344_u0;
reg	[15:0]	syncEnable_u62=16'h0;
reg	[31:0]	syncEnable_u63_u0=32'h0;
reg		reg_6791728c_u0=1'h0;
reg		reg_21434b16_u0=1'h0;
reg	[31:0]	syncEnable_u64_u0=32'h0;
reg	[15:0]	syncEnable_u65_u0=16'h0;
assign add={31'b0, port_3927e736_}+32'h0;
assign and_u1310_u0=reg_21434b16_u0&port_7b58ab67_;
assign subtract={8'b0, port_3927e736_}-9'h1;
assign greaterThanEqualTo_a_signed={subtract[2], subtract[2], subtract[2], subtract[2], subtract[2], subtract[2], subtract[2:0]};
assign greaterThanEqualTo_b_signed=9'h0;
assign greaterThanEqualTo=greaterThanEqualTo_a_signed>=greaterThanEqualTo_b_signed;
assign not_u252_u0=~greaterThanEqualTo;
assign and_u1311_u0=GO&greaterThanEqualTo;
assign and_u1312_u0=GO&not_u252_u0;
assign subtract_u0={8'b0, port_3927e736_}-9'h1;
assign and_u1313_u0=and_u1312_u0&GO;
assign and_u1314_u0=and_u1311_u0&GO;
assign mux_u80=(and_u1314_u0)?{subtract_u0[2], subtract_u0[2], subtract_u0[2], subtract_u0[2], subtract_u0[2], subtract_u0[2], subtract_u0[2:0]}:9'h2;
assign add_u24={mux_u80[2], mux_u80[2], mux_u80[2], mux_u80[2], mux_u80[2], mux_u80[2], mux_u80[2], mux_u80[2], mux_u80[2], mux_u80[2], mux_u80[2], mux_u80[2], mux_u80[2], mux_u80[2], mux_u80[2], mux_u80[2], mux_u80[2], mux_u80[2], mux_u80[2], mux_u80[2], mux_u80[2], mux_u80[2], mux_u80[2], mux_u80[2], mux_u80[2], mux_u80[2], mux_u80[2], mux_u80[2], mux_u80[2], mux_u80[2:0]}+32'h0;
assign and_u1315_u0=reg_21434b16_u0&port_1f3f2d39_;
assign and_u1317_u0=reg_6791728c_u0&port_7b58ab67_;
assign add_u25={syncEnable_u62[15], syncEnable_u62}+{port_129b8bb2_[15], port_129b8bb2_};
assign subtract_u1=syncEnable_u65_u0-add_u25[16:1];
assign simplePinWrite=16'h1&{16{1'h1}};
assign simplePinWrite_u212=subtract_u1&{16{reg_6791728c_u0}};
assign simplePinWrite_u213=reg_6791728c_u0&{1{reg_6791728c_u0}};
assign simplePinWrite_u214=subtract_u1&{16{reg_6791728c_u0}};
assign simplePinWrite_u215=reg_6791728c_u0&{1{reg_6791728c_u0}};
assign simplePinWrite_u216=16'h1&{16{1'h1}};
assign mux_u81_u0=(reg_21434b16_u0)?syncEnable_u63_u0:32'h0;
assign or_u344_u0=reg_21434b16_u0|reg_6791728c_u0;
always @(posedge CLK)
begin
if (reg_21434b16_u0)
syncEnable_u62<=port_1df607d4_;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u63_u0<={add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2:0]};
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6791728c_u0<=1'h0;
else reg_6791728c_u0<=reg_21434b16_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_21434b16_u0<=1'h0;
else reg_21434b16_u0<=GO;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u64_u0<=add_u24;
end
always @(posedge CLK)
begin
if (reg_21434b16_u0)
syncEnable_u65_u0<=port_129b8bb2_;
end
assign RESULT=GO;
assign RESULT_u740=1'h0;
assign RESULT_u741=reg_21434b16_u0;
assign RESULT_u742=syncEnable_u64_u0;
assign RESULT_u743=3'h1;
assign RESULT_u744=or_u344_u0;
assign RESULT_u745=mux_u81_u0;
assign RESULT_u746=3'h1;
assign RESULT_u747=simplePinWrite;
assign RESULT_u748=simplePinWrite_u214;
assign RESULT_u749=simplePinWrite_u213;
assign RESULT_u750=simplePinWrite_u215;
assign RESULT_u751=simplePinWrite_u212;
assign RESULT_u752=simplePinWrite_u216;
assign DONE=reg_6791728c_u0;
endmodule



module image1_iunzip_endianswapper_1edd54fb_(endianswapper_1edd54fb_in, endianswapper_1edd54fb_out);
input	[1:0]	endianswapper_1edd54fb_in;
output	[1:0]	endianswapper_1edd54fb_out;
assign endianswapper_1edd54fb_out=endianswapper_1edd54fb_in;
endmodule



module image1_iunzip_endianswapper_3cf254da_(endianswapper_3cf254da_in, endianswapper_3cf254da_out);
input	[1:0]	endianswapper_3cf254da_in;
output	[1:0]	endianswapper_3cf254da_out;
assign endianswapper_3cf254da_out=endianswapper_3cf254da_in;
endmodule



module image1_iunzip_stateVar_fsmState_image1_iunzip(bus_4c915309_, bus_2d7bb642_, bus_02e4d33b_, bus_3412b614_, bus_0d633a7d_);
input		bus_4c915309_;
input		bus_2d7bb642_;
input		bus_02e4d33b_;
input	[1:0]	bus_3412b614_;
output	[1:0]	bus_0d633a7d_;
wire	[1:0]	endianswapper_1edd54fb_out;
wire	[1:0]	endianswapper_3cf254da_out;
reg	[1:0]	stateVar_fsmState_image1_iunzip_u0=2'h0;
image1_iunzip_endianswapper_1edd54fb_ image1_iunzip_endianswapper_1edd54fb__1(.endianswapper_1edd54fb_in(bus_3412b614_), 
  .endianswapper_1edd54fb_out(endianswapper_1edd54fb_out));
image1_iunzip_endianswapper_3cf254da_ image1_iunzip_endianswapper_3cf254da__1(.endianswapper_3cf254da_in(stateVar_fsmState_image1_iunzip_u0), 
  .endianswapper_3cf254da_out(endianswapper_3cf254da_out));
assign bus_0d633a7d_=endianswapper_3cf254da_out;
always @(posedge bus_4c915309_ or posedge bus_2d7bb642_)
begin
if (bus_2d7bb642_)
stateVar_fsmState_image1_iunzip_u0<=2'h0;
else if (bus_02e4d33b_)
stateVar_fsmState_image1_iunzip_u0<=endianswapper_1edd54fb_out;
end
endmodule



module image1_iunzip_streamFun2(CLK, RESET, GO, port_4da7fcea_, port_5ec353a6_, port_45273060_, port_221c496a_, port_0ebd1361_, port_001ed422_, port_08ebfbc1_, port_587fd1a5_, RESULT, RESULT_u753, RESULT_u754, RESULT_u755, RESULT_u756, RESULT_u757, RESULT_u758, RESULT_u759, RESULT_u760, RESULT_u761, RESULT_u762, RESULT_u763, RESULT_u764, RESULT_u765, RESULT_u766, RESULT_u767, RESULT_u768, RESULT_u769, DONE);
input		CLK;
input		RESET;
input		GO;
input		port_4da7fcea_;
input	[31:0]	port_5ec353a6_;
input		port_45273060_;
input	[15:0]	port_221c496a_;
input		port_0ebd1361_;
input		port_001ed422_;
input	[15:0]	port_08ebfbc1_;
input	[15:0]	port_587fd1a5_;
output		RESULT;
output		RESULT_u753;
output		RESULT_u754;
output	[31:0]	RESULT_u755;
output		RESULT_u756;
output	[31:0]	RESULT_u757;
output	[2:0]	RESULT_u758;
output		RESULT_u759;
output	[31:0]	RESULT_u760;
output	[15:0]	RESULT_u761;
output	[2:0]	RESULT_u762;
output		RESULT_u763;
output	[31:0]	RESULT_u764;
output	[2:0]	RESULT_u765;
output	[15:0]	RESULT_u766;
output		RESULT_u767;
output		RESULT_u768;
output	[15:0]	RESULT_u769;
output		DONE;
wire		simplePinWrite;
wire		and_u1320_u0;
reg		reg_3ae25a28_u0=1'h0;
wire		or_u345_u0;
wire	[31:0]	add;
wire		and_u1321_u0;
wire	[8:0]	subtract;
wire signed	[8:0]	greaterThanEqualTo_a_signed;
wire		greaterThanEqualTo;
wire signed	[8:0]	greaterThanEqualTo_b_signed;
wire		not_u253_u0;
wire		and_u1322_u0;
wire		and_u1323_u0;
wire	[8:0]	subtract_u2;
wire		and_u1324_u0;
wire	[8:0]	mux_u82;
wire		and_u1325_u0;
wire	[31:0]	add_u26;
wire		and_u1326_u0;
wire		and_u1328_u0;
wire	[16:0]	add_u27;
wire	[15:0]	add_u28;
wire	[31:0]	add_u29;
wire		simplePinWrite_u217;
wire	[15:0]	simplePinWrite_u218;
wire	[15:0]	simplePinWrite_u219;
reg	[31:0]	syncEnable_u66=32'h0;
reg	[15:0]	syncEnable_u67_u0=16'h0;
reg	[31:0]	syncEnable_u68_u0=32'h0;
wire	[31:0]	mux_u83_u0;
reg	[15:0]	syncEnable_u69_u0=16'h0;
reg		reg_6adf8b78_u0=1'h0;
wire	[31:0]	mux_u84_u0;
wire		or_u346_u0;
reg	[15:0]	syncEnable_u70_u0=16'h0;
reg		reg_26b6f167_u0=1'h0;
reg		reg_26b6f167_result_delayed_u0=1'h0;
assign simplePinWrite=GO&{1{GO}};
assign and_u1320_u0=reg_3ae25a28_u0&port_0ebd1361_;
always @(posedge CLK or posedge reg_26b6f167_u0 or posedge or_u345_u0)
begin
if (or_u345_u0)
reg_3ae25a28_u0<=1'h0;
else if (reg_26b6f167_u0)
reg_3ae25a28_u0<=1'h1;
else reg_3ae25a28_u0<=reg_3ae25a28_u0;
end
assign or_u345_u0=and_u1320_u0|RESET;
assign add={31'b0, port_4da7fcea_}+32'h0;
assign and_u1321_u0=reg_26b6f167_result_delayed_u0&port_001ed422_;
assign subtract={8'b0, port_4da7fcea_}-9'h1;
assign greaterThanEqualTo_a_signed={subtract[2], subtract[2], subtract[2], subtract[2], subtract[2], subtract[2], subtract[2:0]};
assign greaterThanEqualTo_b_signed=9'h0;
assign greaterThanEqualTo=greaterThanEqualTo_a_signed>=greaterThanEqualTo_b_signed;
assign not_u253_u0=~greaterThanEqualTo;
assign and_u1322_u0=GO&greaterThanEqualTo;
assign and_u1323_u0=GO&not_u253_u0;
assign subtract_u2={8'b0, port_4da7fcea_}-9'h1;
assign and_u1324_u0=and_u1323_u0&GO;
assign mux_u82=(and_u1324_u0)?9'h2:{subtract_u2[2], subtract_u2[2], subtract_u2[2], subtract_u2[2], subtract_u2[2], subtract_u2[2], subtract_u2[2:0]};
assign and_u1325_u0=and_u1322_u0&GO;
assign add_u26={mux_u82[2], mux_u82[2], mux_u82[2], mux_u82[2], mux_u82[2], mux_u82[2], mux_u82[2], mux_u82[2], mux_u82[2], mux_u82[2], mux_u82[2], mux_u82[2], mux_u82[2], mux_u82[2], mux_u82[2], mux_u82[2], mux_u82[2], mux_u82[2], mux_u82[2], mux_u82[2], mux_u82[2], mux_u82[2], mux_u82[2], mux_u82[2], mux_u82[2], mux_u82[2], mux_u82[2], mux_u82[2], mux_u82[2], mux_u82[2:0]}+32'h0;
assign and_u1326_u0=reg_26b6f167_result_delayed_u0&port_0ebd1361_;
assign and_u1328_u0=reg_6adf8b78_u0&port_001ed422_;
assign add_u27={syncEnable_u67_u0[15], syncEnable_u67_u0}+{port_08ebfbc1_[15], port_08ebfbc1_};
assign add_u28=syncEnable_u69_u0+{add_u27[16], add_u27[16:2]};
assign add_u29=port_5ec353a6_+32'h1;
assign simplePinWrite_u217=reg_6adf8b78_u0&{1{reg_6adf8b78_u0}};
assign simplePinWrite_u218=16'h1&{16{1'h1}};
assign simplePinWrite_u219=add_u28&{16{reg_6adf8b78_u0}};
always @(posedge CLK)
begin
if (GO)
syncEnable_u66<={add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2:0]};
end
always @(posedge CLK)
begin
if (reg_26b6f167_result_delayed_u0)
syncEnable_u67_u0<=port_221c496a_;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u68_u0<=add_u26;
end
assign mux_u83_u0=(reg_26b6f167_u0)?32'h0:syncEnable_u68_u0;
always @(posedge CLK)
begin
if (reg_26b6f167_result_delayed_u0)
syncEnable_u69_u0<=port_08ebfbc1_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6adf8b78_u0<=1'h0;
else reg_6adf8b78_u0<=reg_26b6f167_result_delayed_u0;
end
assign mux_u84_u0=(reg_26b6f167_result_delayed_u0)?syncEnable_u66:32'h0;
assign or_u346_u0=reg_26b6f167_result_delayed_u0|reg_6adf8b78_u0;
always @(posedge CLK)
begin
if (GO)
syncEnable_u70_u0<=port_587fd1a5_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_26b6f167_u0<=1'h0;
else reg_26b6f167_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_26b6f167_result_delayed_u0<=1'h0;
else reg_26b6f167_result_delayed_u0<=reg_26b6f167_u0;
end
assign RESULT=GO;
assign RESULT_u753=1'h0;
assign RESULT_u754=GO;
assign RESULT_u755=add_u29;
assign RESULT_u756=reg_26b6f167_result_delayed_u0;
assign RESULT_u757=mux_u83_u0;
assign RESULT_u758=3'h1;
assign RESULT_u759=reg_26b6f167_u0;
assign RESULT_u760=mux_u83_u0;
assign RESULT_u761=syncEnable_u70_u0;
assign RESULT_u762=3'h1;
assign RESULT_u763=or_u346_u0;
assign RESULT_u764=mux_u84_u0;
assign RESULT_u765=3'h1;
assign RESULT_u766=simplePinWrite_u219;
assign RESULT_u767=simplePinWrite_u217;
assign RESULT_u768=simplePinWrite;
assign RESULT_u769=simplePinWrite_u218;
assign DONE=reg_6adf8b78_u0;
endmodule



module image1_iunzip_stateVar_midPoint(bus_676a86b4_, bus_7f9b1e16_, bus_6d113f7e_, bus_79b19529_, bus_196aa05d_, bus_5894ff4e_, bus_4ddfe8ac_, bus_56ab03e3_, bus_3b63cd45_, bus_4ba5b0a8_, bus_79302887_);
input		bus_676a86b4_;
input		bus_7f9b1e16_;
input		bus_6d113f7e_;
input		bus_79b19529_;
input		bus_196aa05d_;
input		bus_5894ff4e_;
input		bus_4ddfe8ac_;
input		bus_56ab03e3_;
input		bus_3b63cd45_;
input		bus_4ba5b0a8_;
output		bus_79302887_;
wire		or_29667c9f_u0;
reg		stateVar_midPoint_u0=1'h1;
assign bus_79302887_=stateVar_midPoint_u0;
assign or_29667c9f_u0=bus_6d113f7e_|bus_196aa05d_|bus_4ddfe8ac_|bus_3b63cd45_;
always @(posedge bus_676a86b4_ or posedge bus_7f9b1e16_)
begin
if (bus_7f9b1e16_)
stateVar_midPoint_u0<=1'h1;
else if (or_29667c9f_u0)
stateVar_midPoint_u0<=1'h0;
end
endmodule



module image1_iunzip_endianswapper_70c883ac_(endianswapper_70c883ac_in, endianswapper_70c883ac_out);
input	[31:0]	endianswapper_70c883ac_in;
output	[31:0]	endianswapper_70c883ac_out;
assign endianswapper_70c883ac_out=endianswapper_70c883ac_in;
endmodule



module image1_iunzip_endianswapper_3e51e7fe_(endianswapper_3e51e7fe_in, endianswapper_3e51e7fe_out);
input	[31:0]	endianswapper_3e51e7fe_in;
output	[31:0]	endianswapper_3e51e7fe_out;
assign endianswapper_3e51e7fe_out=endianswapper_3e51e7fe_in;
endmodule



module image1_iunzip_stateVar_In1TokenIndex(bus_00a6f1a7_, bus_05ce656d_, bus_69335eb2_, bus_28bc525f_, bus_6bbd8c15_);
input		bus_00a6f1a7_;
input		bus_05ce656d_;
input		bus_69335eb2_;
input	[31:0]	bus_28bc525f_;
output	[31:0]	bus_6bbd8c15_;
wire	[31:0]	endianswapper_70c883ac_out;
reg	[31:0]	stateVar_In1TokenIndex_u0=32'h0;
wire	[31:0]	endianswapper_3e51e7fe_out;
image1_iunzip_endianswapper_70c883ac_ image1_iunzip_endianswapper_70c883ac__1(.endianswapper_70c883ac_in(bus_28bc525f_), 
  .endianswapper_70c883ac_out(endianswapper_70c883ac_out));
assign bus_6bbd8c15_=endianswapper_3e51e7fe_out;
always @(posedge bus_00a6f1a7_ or posedge bus_05ce656d_)
begin
if (bus_05ce656d_)
stateVar_In1TokenIndex_u0<=32'h0;
else if (bus_69335eb2_)
stateVar_In1TokenIndex_u0<=endianswapper_70c883ac_out;
end
image1_iunzip_endianswapper_3e51e7fe_ image1_iunzip_endianswapper_3e51e7fe__1(.endianswapper_3e51e7fe_in(stateVar_In1TokenIndex_u0), 
  .endianswapper_3e51e7fe_out(endianswapper_3e51e7fe_out));
endmodule



module image1_iunzip_endianswapper_01b25bf2_(endianswapper_01b25bf2_in, endianswapper_01b25bf2_out);
input	[31:0]	endianswapper_01b25bf2_in;
output	[31:0]	endianswapper_01b25bf2_out;
assign endianswapper_01b25bf2_out={endianswapper_01b25bf2_in[31:2], 1'b1, endianswapper_01b25bf2_in[0]};
endmodule



module image1_iunzip_endianswapper_0f9a6f77_(endianswapper_0f9a6f77_in, endianswapper_0f9a6f77_out);
input	[31:0]	endianswapper_0f9a6f77_in;
output	[31:0]	endianswapper_0f9a6f77_out;
assign endianswapper_0f9a6f77_out=endianswapper_0f9a6f77_in;
endmodule



module image1_iunzip_stateVar_In1MaxTokenIndex(bus_022df17c_, bus_1facd4e4_, bus_4a9eda6d_, bus_5e278fb9_, bus_6d8ec6c0_);
input		bus_022df17c_;
input		bus_1facd4e4_;
input		bus_4a9eda6d_;
input	[31:0]	bus_5e278fb9_;
output	[31:0]	bus_6d8ec6c0_;
wire	[31:0]	endianswapper_01b25bf2_out;
reg	[31:0]	stateVar_In1MaxTokenIndex_u0=32'h0;
wire	[31:0]	endianswapper_0f9a6f77_out;
image1_iunzip_endianswapper_01b25bf2_ image1_iunzip_endianswapper_01b25bf2__1(.endianswapper_01b25bf2_in({bus_5e278fb9_[31:2], 1'b0, bus_5e278fb9_[0]}), 
  .endianswapper_01b25bf2_out(endianswapper_01b25bf2_out));
assign bus_6d8ec6c0_=endianswapper_0f9a6f77_out;
always @(posedge bus_022df17c_ or posedge bus_1facd4e4_)
begin
if (bus_1facd4e4_)
stateVar_In1MaxTokenIndex_u0<=32'h0;
else if (bus_4a9eda6d_)
stateVar_In1MaxTokenIndex_u0<={endianswapper_01b25bf2_out[31:2], 1'b1, endianswapper_01b25bf2_out[0]};
end
image1_iunzip_endianswapper_0f9a6f77_ image1_iunzip_endianswapper_0f9a6f77__1(.endianswapper_0f9a6f77_in(stateVar_In1MaxTokenIndex_u0), 
  .endianswapper_0f9a6f77_out(endianswapper_0f9a6f77_out));
endmodule



module image1_iunzip_simplememoryreferee_0b0f52d7_(bus_29cdd1f8_, bus_6b72c155_, bus_3c855b7b_, bus_20f0729f_, bus_5b77758f_, bus_5b45fa2c_, bus_0964b8c9_, bus_37539c61_, bus_1daba9ee_, bus_0e50a633_, bus_6d9883cb_, bus_5525d2cf_, bus_5038a20c_, bus_267b146b_, bus_67995a05_, bus_5fbad179_, bus_5f260ad4_, bus_711ba866_, bus_3d439865_, bus_2e00db39_, bus_3f0f2b61_, bus_1de509a3_, bus_438eba07_, bus_01bb560e_, bus_3c8caa47_, bus_349fc2ad_, bus_7818c025_, bus_185cf169_, bus_380af87e_);
input		bus_29cdd1f8_;
input		bus_6b72c155_;
input		bus_3c855b7b_;
input	[15:0]	bus_20f0729f_;
input		bus_5b77758f_;
input	[31:0]	bus_5b45fa2c_;
input	[2:0]	bus_0964b8c9_;
input		bus_37539c61_;
input	[31:0]	bus_1daba9ee_;
input	[2:0]	bus_0e50a633_;
input		bus_6d9883cb_;
input	[31:0]	bus_5525d2cf_;
input	[2:0]	bus_5038a20c_;
input		bus_267b146b_;
input	[31:0]	bus_67995a05_;
input	[2:0]	bus_5fbad179_;
output	[15:0]	bus_5f260ad4_;
output	[31:0]	bus_711ba866_;
output		bus_3d439865_;
output		bus_2e00db39_;
output	[2:0]	bus_3f0f2b61_;
output	[15:0]	bus_1de509a3_;
output		bus_438eba07_;
output	[15:0]	bus_01bb560e_;
output		bus_3c8caa47_;
output	[15:0]	bus_349fc2ad_;
output		bus_7818c025_;
output	[15:0]	bus_185cf169_;
output		bus_380af87e_;
wire		or_713ef07e_u0;
reg		done_qual_u42=1'h0;
wire		and_72584599_u0;
wire		or_27a047aa_u0;
wire		or_45f26528_u0;
wire		not_029b83c1_u0;
wire		and_08cc2292_u0;
wire		and_6d00581f_u0;
wire		not_03e44387_u0;
reg		done_qual_u43_u0=1'h0;
reg		done_qual_u44_u0=1'h0;
wire		or_38b1f2dd_u0;
wire		and_53170f7a_u0;
wire		not_6cc0952e_u0;
reg		done_qual_u45_u0=1'h0;
wire		not_7be34452_u0;
wire	[31:0]	mux_5016beae_u0;
wire		or_7734ba4e_u0;
assign or_713ef07e_u0=bus_5b77758f_|bus_37539c61_|bus_6d9883cb_|bus_267b146b_;
always @(posedge bus_29cdd1f8_)
begin
if (bus_6b72c155_)
done_qual_u42<=1'h0;
else done_qual_u42<=bus_5b77758f_;
end
assign and_72584599_u0=or_7734ba4e_u0&bus_3c855b7b_;
assign or_27a047aa_u0=bus_37539c61_|done_qual_u43_u0;
assign or_45f26528_u0=bus_5b77758f_|done_qual_u42;
assign not_029b83c1_u0=~bus_3c855b7b_;
assign and_08cc2292_u0=or_27a047aa_u0&bus_3c855b7b_;
assign and_6d00581f_u0=or_45f26528_u0&bus_3c855b7b_;
assign not_03e44387_u0=~bus_3c855b7b_;
always @(posedge bus_29cdd1f8_)
begin
if (bus_6b72c155_)
done_qual_u43_u0<=1'h0;
else done_qual_u43_u0<=bus_37539c61_;
end
assign bus_5f260ad4_=16'h0;
assign bus_711ba866_=mux_5016beae_u0;
assign bus_3d439865_=1'h0;
assign bus_2e00db39_=or_713ef07e_u0;
assign bus_3f0f2b61_=3'h1;
assign bus_1de509a3_=bus_20f0729f_;
assign bus_438eba07_=and_6d00581f_u0;
assign bus_01bb560e_=bus_20f0729f_;
assign bus_3c8caa47_=and_08cc2292_u0;
assign bus_349fc2ad_=bus_20f0729f_;
assign bus_7818c025_=and_53170f7a_u0;
assign bus_185cf169_=bus_20f0729f_;
assign bus_380af87e_=and_72584599_u0;
always @(posedge bus_29cdd1f8_)
begin
if (bus_6b72c155_)
done_qual_u44_u0<=1'h0;
else done_qual_u44_u0<=bus_6d9883cb_;
end
assign or_38b1f2dd_u0=bus_6d9883cb_|done_qual_u44_u0;
assign and_53170f7a_u0=or_38b1f2dd_u0&bus_3c855b7b_;
assign not_6cc0952e_u0=~bus_3c855b7b_;
always @(posedge bus_29cdd1f8_)
begin
if (bus_6b72c155_)
done_qual_u45_u0<=1'h0;
else done_qual_u45_u0<=bus_267b146b_;
end
assign not_7be34452_u0=~bus_3c855b7b_;
assign mux_5016beae_u0=({32{bus_5b77758f_}}&bus_5b45fa2c_)|({32{bus_37539c61_}}&bus_1daba9ee_)|({32{bus_6d9883cb_}}&bus_5525d2cf_)|({32{bus_267b146b_}}&bus_67995a05_);
assign or_7734ba4e_u0=bus_267b146b_|done_qual_u45_u0;
endmodule



module image1_iunzip_streamFun1(CLK, RESET, GO, port_4691c47d_, port_0289ded9_, port_635f8008_, port_747b457f_, port_1d854cce_, port_7ab2bf13_, port_6ecc5cde_, port_01e6d96a_, RESULT, RESULT_u770, RESULT_u771, RESULT_u772, RESULT_u773, RESULT_u774, RESULT_u775, RESULT_u776, RESULT_u777, RESULT_u778, RESULT_u779, RESULT_u780, RESULT_u781, RESULT_u782, RESULT_u783, RESULT_u784, RESULT_u785, RESULT_u786, DONE);
input		CLK;
input		RESET;
input		GO;
input		port_4691c47d_;
input	[31:0]	port_0289ded9_;
input		port_635f8008_;
input	[15:0]	port_747b457f_;
input		port_1d854cce_;
input		port_7ab2bf13_;
input	[15:0]	port_6ecc5cde_;
input	[15:0]	port_01e6d96a_;
output		RESULT;
output		RESULT_u770;
output		RESULT_u771;
output	[31:0]	RESULT_u772;
output		RESULT_u773;
output	[31:0]	RESULT_u774;
output	[2:0]	RESULT_u775;
output		RESULT_u776;
output	[31:0]	RESULT_u777;
output	[15:0]	RESULT_u778;
output	[2:0]	RESULT_u779;
output		RESULT_u780;
output	[31:0]	RESULT_u781;
output	[2:0]	RESULT_u782;
output	[15:0]	RESULT_u783;
output		RESULT_u784;
output	[15:0]	RESULT_u785;
output		RESULT_u786;
output		DONE;
wire		simplePinWrite;
wire		or_u347_u0;
wire		and_u1331_u0;
reg		reg_55d15bea_u0=1'h0;
wire	[31:0]	add;
wire		and_u1332_u0;
wire	[8:0]	subtract;
wire signed	[8:0]	greaterThanEqualTo_a_signed;
wire		greaterThanEqualTo;
wire signed	[8:0]	greaterThanEqualTo_b_signed;
wire		not_u254_u0;
wire		and_u1333_u0;
wire		and_u1334_u0;
wire	[8:0]	subtract_u3;
wire		and_u1335_u0;
wire		and_u1336_u0;
wire	[8:0]	mux_u85;
wire	[31:0]	add_u30;
wire		and_u1337_u0;
wire		and_u1339_u0;
wire	[16:0]	add_u31;
wire	[15:0]	subtract_u4;
wire	[31:0]	add_u32;
wire		simplePinWrite_u220;
wire	[15:0]	simplePinWrite_u221;
wire	[15:0]	simplePinWrite_u222;
wire	[31:0]	mux_u86_u0;
wire		or_u348_u0;
reg		reg_2aa4b998_u0=1'h0;
reg	[31:0]	syncEnable_u71=32'h0;
reg	[15:0]	syncEnable_u72_u0=16'h0;
reg	[15:0]	syncEnable_u73_u0=16'h0;
reg	[31:0]	syncEnable_u74_u0=32'h0;
reg		reg_4b98de26_u0=1'h0;
reg	[15:0]	syncEnable_u75_u0=16'h0;
wire	[31:0]	mux_u87_u0;
reg		reg_4b98de26_result_delayed_u0=1'h0;
assign simplePinWrite=GO&{1{GO}};
assign or_u347_u0=and_u1331_u0|RESET;
assign and_u1331_u0=reg_55d15bea_u0&port_1d854cce_;
always @(posedge CLK or posedge reg_4b98de26_u0 or posedge or_u347_u0)
begin
if (or_u347_u0)
reg_55d15bea_u0<=1'h0;
else if (reg_4b98de26_u0)
reg_55d15bea_u0<=1'h1;
else reg_55d15bea_u0<=reg_55d15bea_u0;
end
assign add={31'b0, port_4691c47d_}+32'h0;
assign and_u1332_u0=reg_4b98de26_result_delayed_u0&port_7ab2bf13_;
assign subtract={8'b0, port_4691c47d_}-9'h1;
assign greaterThanEqualTo_a_signed={subtract[2], subtract[2], subtract[2], subtract[2], subtract[2], subtract[2], subtract[2:0]};
assign greaterThanEqualTo_b_signed=9'h0;
assign greaterThanEqualTo=greaterThanEqualTo_a_signed>=greaterThanEqualTo_b_signed;
assign not_u254_u0=~greaterThanEqualTo;
assign and_u1333_u0=GO&greaterThanEqualTo;
assign and_u1334_u0=GO&not_u254_u0;
assign subtract_u3={8'b0, port_4691c47d_}-9'h1;
assign and_u1335_u0=and_u1333_u0&GO;
assign and_u1336_u0=and_u1334_u0&GO;
assign mux_u85=(and_u1336_u0)?9'h2:{subtract_u3[2], subtract_u3[2], subtract_u3[2], subtract_u3[2], subtract_u3[2], subtract_u3[2], subtract_u3[2:0]};
assign add_u30={mux_u85[2], mux_u85[2], mux_u85[2], mux_u85[2], mux_u85[2], mux_u85[2], mux_u85[2], mux_u85[2], mux_u85[2], mux_u85[2], mux_u85[2], mux_u85[2], mux_u85[2], mux_u85[2], mux_u85[2], mux_u85[2], mux_u85[2], mux_u85[2], mux_u85[2], mux_u85[2], mux_u85[2], mux_u85[2], mux_u85[2], mux_u85[2], mux_u85[2], mux_u85[2], mux_u85[2], mux_u85[2], mux_u85[2], mux_u85[2:0]}+32'h0;
assign and_u1337_u0=reg_4b98de26_result_delayed_u0&port_1d854cce_;
assign and_u1339_u0=reg_2aa4b998_u0&port_7ab2bf13_;
assign add_u31={syncEnable_u73_u0[15], syncEnable_u73_u0}+{port_6ecc5cde_[15], port_6ecc5cde_};
assign subtract_u4=syncEnable_u72_u0-add_u31[16:1];
assign add_u32=port_0289ded9_+32'h1;
assign simplePinWrite_u220=reg_2aa4b998_u0&{1{reg_2aa4b998_u0}};
assign simplePinWrite_u221=subtract_u4&{16{reg_2aa4b998_u0}};
assign simplePinWrite_u222=16'h1&{16{1'h1}};
assign mux_u86_u0=(reg_4b98de26_result_delayed_u0)?syncEnable_u74_u0:32'h0;
assign or_u348_u0=reg_4b98de26_result_delayed_u0|reg_2aa4b998_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2aa4b998_u0<=1'h0;
else reg_2aa4b998_u0<=reg_4b98de26_result_delayed_u0;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u71<=add_u30;
end
always @(posedge CLK)
begin
if (reg_4b98de26_result_delayed_u0)
syncEnable_u72_u0<=port_6ecc5cde_;
end
always @(posedge CLK)
begin
if (reg_4b98de26_result_delayed_u0)
syncEnable_u73_u0<=port_747b457f_;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u74_u0<={add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2:0]};
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4b98de26_u0<=1'h0;
else reg_4b98de26_u0<=GO;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u75_u0<=port_01e6d96a_;
end
assign mux_u87_u0=(reg_4b98de26_u0)?32'h0:syncEnable_u71;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4b98de26_result_delayed_u0<=1'h0;
else reg_4b98de26_result_delayed_u0<=reg_4b98de26_u0;
end
assign RESULT=GO;
assign RESULT_u770=1'h0;
assign RESULT_u771=GO;
assign RESULT_u772=add_u32;
assign RESULT_u773=reg_4b98de26_result_delayed_u0;
assign RESULT_u774=mux_u87_u0;
assign RESULT_u775=3'h1;
assign RESULT_u776=reg_4b98de26_u0;
assign RESULT_u777=mux_u87_u0;
assign RESULT_u778=syncEnable_u75_u0;
assign RESULT_u779=3'h1;
assign RESULT_u780=or_u348_u0;
assign RESULT_u781=mux_u86_u0;
assign RESULT_u782=3'h1;
assign RESULT_u783=simplePinWrite_u222;
assign RESULT_u784=simplePinWrite_u220;
assign RESULT_u785=simplePinWrite_u221;
assign RESULT_u786=simplePinWrite;
assign DONE=reg_2aa4b998_u0;
endmodule



module image1_iunzip_simplememoryreferee_4f4a8814_(bus_6a794fd6_, bus_561f7191_, bus_495872da_, bus_220964f4_, bus_31862682_, bus_0040cf15_, bus_5ccabeca_, bus_56d7b0af_, bus_59b1b34a_, bus_5b4fce35_, bus_4d510363_, bus_6aac9d02_, bus_3f4ce93d_, bus_4ef7394f_);
input		bus_6a794fd6_;
input		bus_561f7191_;
input		bus_495872da_;
input	[15:0]	bus_220964f4_;
input		bus_31862682_;
input	[31:0]	bus_0040cf15_;
input	[2:0]	bus_5ccabeca_;
output	[15:0]	bus_56d7b0af_;
output	[31:0]	bus_59b1b34a_;
output		bus_5b4fce35_;
output		bus_4d510363_;
output	[2:0]	bus_6aac9d02_;
output	[15:0]	bus_3f4ce93d_;
output		bus_4ef7394f_;
assign bus_56d7b0af_=16'h0;
assign bus_59b1b34a_=32'h1;
assign bus_5b4fce35_=1'h0;
assign bus_4d510363_=bus_31862682_;
assign bus_6aac9d02_=3'h1;
assign bus_3f4ce93d_=bus_220964f4_;
assign bus_4ef7394f_=bus_495872da_;
endmodule



module image1_iunzip_Kicker_22(CLK, RESET, bus_0532da99_);
input		CLK;
input		RESET;
output		bus_0532da99_;
wire		bus_23009074_;
reg		kicker_1=1'h0;
reg		kicker_res=1'h0;
wire		bus_3884fe31_;
wire		bus_1ec24681_;
reg		kicker_2=1'h0;
wire		bus_6d7766e3_;
assign bus_23009074_=~kicker_2;
always @(posedge CLK)
begin
kicker_1<=bus_6d7766e3_;
end
always @(posedge CLK)
begin
kicker_res<=bus_3884fe31_;
end
assign bus_3884fe31_=kicker_1&bus_6d7766e3_&bus_23009074_;
assign bus_1ec24681_=bus_6d7766e3_&kicker_1;
always @(posedge CLK)
begin
kicker_2<=bus_1ec24681_;
end
assign bus_0532da99_=kicker_res;
assign bus_6d7766e3_=~RESET;
endmodule



module image1_iunzip_scheduler(CLK, RESET, GO, port_18e00d02_, port_7b9868d2_, port_5b5cde36_, port_7a3e2d5e_, port_2b235147_, port_30bf0bb1_, port_2d451d49_, port_01ffd1e5_, port_6c59504e_, port_7dc7ca1e_, port_2f06a0cc_, port_2cc0cc2a_, port_65a60be6_, port_0312d0b7_, port_4fbbb17b_, RESULT, RESULT_u787, RESULT_u788, RESULT_u789, RESULT_u790, RESULT_u791, RESULT_u792, RESULT_u793, RESULT_u794, RESULT_u795, RESULT_u796, RESULT_u797, RESULT_u798, RESULT_u799, RESULT_u800, RESULT_u801, RESULT_u802, RESULT_u803, RESULT_u804, RESULT_u805, DONE);
input		CLK;
input		RESET;
input		GO;
input	[1:0]	port_18e00d02_;
input	[1:0]	port_7b9868d2_;
input	[31:0]	port_5b5cde36_;
input	[31:0]	port_7a3e2d5e_;
input	[31:0]	port_2b235147_;
input		port_30bf0bb1_;
input		port_2d451d49_;
input		port_01ffd1e5_;
input		port_6c59504e_;
input	[15:0]	port_7dc7ca1e_;
input		port_2f06a0cc_;
input		port_2cc0cc2a_;
input		port_65a60be6_;
input		port_0312d0b7_;
input		port_4fbbb17b_;
output		RESULT;
output	[1:0]	RESULT_u787;
output		RESULT_u788;
output	[1:0]	RESULT_u789;
output		RESULT_u790;
output	[31:0]	RESULT_u791;
output		RESULT_u792;
output	[31:0]	RESULT_u793;
output		RESULT_u794;
output		RESULT_u795;
output		RESULT_u796;
output	[31:0]	RESULT_u797;
output	[15:0]	RESULT_u798;
output	[2:0]	RESULT_u799;
output		RESULT_u800;
output		RESULT_u801;
output		RESULT_u802;
output		RESULT_u803;
output		RESULT_u804;
output		RESULT_u805;
output		DONE;
wire		and_u1341_u0;
wire signed	[31:0]	equals_a_signed;
wire signed	[31:0]	equals_b_signed;
wire		equals;
wire		equals_u74;
wire signed	[31:0]	equals_u74_b_signed;
wire signed	[31:0]	equals_u74_a_signed;
wire signed	[31:0]	equals_u75_b_signed;
wire		equals_u75;
wire signed	[31:0]	equals_u75_a_signed;
wire signed	[31:0]	equals_u76_b_signed;
wire		equals_u76;
wire signed	[31:0]	equals_u76_a_signed;
wire		and_u1342_u0;
wire		and_u1343_u0;
wire		not_u255_u0;
wire		and_u1344_u0;
wire		not_u256_u0;
wire		and_u1345_u0;
wire		simplePinWrite;
reg		reg_55828783_u0=1'h0;
reg		reg_39bf2b99_u0=1'h0;
reg		reg_39bf2b99_result_delayed_u0=1'h0;
wire		and_u1346_u0;
wire		or_u349_u0;
reg		reg_39bf2b99_result_delayed_result_delayed_u0=1'h0;
wire		and_u1347_u0;
wire	[1:0]	mux_u88;
wire		or_u350_u0;
wire		or_u351_u0;
wire		and_u1348_u0;
reg		and_delayed_u71=1'h0;
wire		and_u1349_u0;
wire signed	[31:0]	equals_u77_a_signed;
wire		equals_u77;
wire signed	[31:0]	equals_u77_b_signed;
wire		not_u257_u0;
wire		and_u1350_u0;
wire		and_u1351_u0;
wire		and_u1352_u0;
wire		and_u1353_u0;
wire		not_u258_u0;
wire		andOp;
wire		not_u259_u0;
wire		and_u1354_u0;
wire		and_u1355_u0;
wire		simplePinWrite_u223;
wire		or_u352_u0;
wire		and_u1356_u0;
reg		reg_49e39485_u0=1'h0;
reg		and_delayed_u72_u0=1'h0;
wire		and_u1357_u0;
reg		and_delayed_u73_u0=1'h0;
wire		and_u1358_u0;
wire		not_u260_u0;
wire		and_u1359_u0;
wire		and_u1360_u0;
wire		not_u261_u0;
wire		and_u1361_u0;
wire		simplePinWrite_u224;
wire		or_u353_u0;
reg		reg_7a1ee0d6_u0=1'h0;
wire		and_u1362_u0;
reg		reg_7bb2e7de_u0=1'h0;
reg		reg_64307160_u0=1'h0;
wire		and_u1363_u0;
reg		and_delayed_u74_u0=1'h0;
wire		and_u1364_u0;
wire		or_u354_u0;
wire		and_u1365_u0;
reg		and_delayed_u75_u0=1'h0;
wire	[1:0]	mux_u89_u0;
wire		or_u355_u0;
wire		or_u356_u0;
wire	[1:0]	mux_u90_u0;
wire		or_u357_u0;
wire		and_u1366_u0;
wire		and_u1367_u0;
reg		reg_00382bbc_u0=1'h0;
wire		and_u1368_u0;
wire		or_u358_u0;
wire		and_u1369_u0;
wire		equals_u78;
wire signed	[31:0]	equals_u78_a_signed;
wire signed	[31:0]	equals_u78_b_signed;
wire		and_u1370_u0;
wire		and_u1371_u0;
wire		not_u262_u0;
wire		and_u1372_u0;
wire		not_u263_u0;
wire		and_u1373_u0;
wire		andOp_u108;
wire		and_u1374_u0;
wire		not_u264_u0;
wire		and_u1375_u0;
wire		simplePinWrite_u225;
wire		and_u1376_u0;
wire		and_u1377_u0;
reg		reg_04ddc90f_u0=1'h0;
reg		and_delayed_u76_u0=1'h0;
wire		or_u359_u0;
reg		and_delayed_u77_u0=1'h0;
wire		not_u265_u0;
wire		and_u1378_u0;
wire		and_u1379_u0;
wire		and_u1380_u0;
wire		not_u266_u0;
wire		and_u1381_u0;
wire		simplePinWrite_u226;
reg		reg_5ed9e738_u0=1'h0;
reg		reg_679f5f5d_u0=1'h0;
wire		or_u360_u0;
reg		reg_5ed9e738_result_delayed_u0=1'h0;
wire		and_u1382_u0;
wire		and_u1383_u0;
reg		and_delayed_u78_u0=1'h0;
reg		reg_5cab12fe_u0=1'h0;
wire		and_u1384_u0;
wire		or_u361_u0;
wire	[1:0]	mux_u91_u0;
wire		or_u362_u0;
wire		and_u1385_u0;
wire		and_u1386_u0;
wire		and_u1387_u0;
wire		or_u363_u0;
wire		or_u364_u0;
wire	[1:0]	mux_u92_u0;
reg		reg_29f791b4_u0=1'h0;
wire		and_u1388_u0;
wire		or_u365_u0;
wire		and_u1389_u0;
wire signed	[31:0]	equals_u79_b_signed;
wire		equals_u79;
wire signed	[31:0]	equals_u79_a_signed;
wire		and_u1390_u0;
wire		and_u1391_u0;
wire		not_u267_u0;
wire signed	[31:0]	lessThan_b_signed;
wire signed	[31:0]	lessThan_a_signed;
wire		lessThan;
wire		not_u268_u0;
wire		and_u1392_u0;
wire		and_u1393_u0;
wire		and_u1394_u0;
wire		not_u269_u0;
wire		and_u1395_u0;
wire		simplePinWrite_u227;
wire	[31:0]	add;
reg		reg_22328357_u0=1'h0;
wire		or_u366_u0;
wire		and_u1396_u0;
wire	[31:0]	add_u33;
reg	[15:0]	syncEnable_u76=16'h0;
wire		and_u1397_u0;
wire	[15:0]	mux_u93_u0;
wire		and_u1398_u0;
reg	[15:0]	syncEnable_u77_u0=16'h0;
reg		and_delayed_u79_u0=1'h0;
reg		and_delayed_u80_u0=1'h0;
reg	[2:0]	syncEnable_u78_u0=3'h0;
reg	[15:0]	syncEnable_u79_u0=16'h0;
wire		and_u1399_u0;
wire	[15:0]	mux_u94_u0;
reg	[31:0]	syncEnable_u80_u0=32'h0;
wire		and_u1400_u0;
reg		and_delayed_u81_u0=1'h0;
reg		and_delayed_u82_u0=1'h0;
wire	[31:0]	mux_u95_u0;
wire	[15:0]	mux_u96_u0;
wire	[31:0]	mux_u97_u0;
wire		and_u1401_u0;
wire		and_u1402_u0;
reg		and_delayed_u83_u0=1'h0;
reg		and_delayed_u84_u0=1'h0;
reg	[15:0]	syncEnable_u81_u0=16'h0;
reg	[31:0]	syncEnable_u82_u0=32'h0;
wire	[31:0]	latch_1f7403f6_out;
reg	[31:0]	latch_1f7403f6_reg=32'h0;
wire		or_u367_u0;
wire	[31:0]	mux_u98_u0;
wire		or_u368_u0;
wire	[1:0]	mux_u99_u0;
wire	[1:0]	mux_u100_u0;
wire		or_u369_u0;
wire		or_u370_u0;
wire	[31:0]	mux_u101_u0;
reg		scoreboard_428a1a5c_reg1=1'h0;
wire		scoreboard_428a1a5c_resOr0;
wire		scoreboard_428a1a5c_and;
wire		scoreboard_428a1a5c_resOr1;
wire		bus_3c51dea1_;
reg		scoreboard_428a1a5c_reg0=1'h0;
reg		scoreboard_428a1a5c_reg2=1'h0;
wire		scoreboard_428a1a5c_resOr2;
reg	[15:0]	latch_7da74311_reg=16'h0;
wire	[15:0]	latch_7da74311_out;
reg		block_GO_delayed_u0=1'h0;
reg		syncEnable_u83_u0=1'h0;
reg		syncEnable_u84_u0=1'h0;
reg		syncEnable_u85_u0=1'h0;
reg	[31:0]	syncEnable_u86_u0=32'h0;
reg	[31:0]	syncEnable_u87_u0=32'h0;
reg		syncEnable_u88_u0=1'h0;
reg	[2:0]	syncEnable_u89_u0=3'h0;
reg		syncEnable_u90_u0=1'h0;
reg	[31:0]	syncEnable_u91_u0=32'h0;
reg		syncEnable_u92_u0=1'h0;
reg	[15:0]	syncEnable_u93_u0=16'h0;
reg		block_GO_delayed_u1_u0=1'h0;
wire	[15:0]	mux_u102_u0;
reg	[31:0]	fbReg_temp_fsmOldState_image1_iunzip_0_u0=32'h0;
reg	[15:0]	fbReg_In1Portvalue_u0=16'h0;
reg		syncEnable_u94_u0=1'h0;
reg		loopControl_u0=1'h0;
wire		or_u371_u0;
wire	[31:0]	mux_u103_u0;
reg		reg_65426ec1_u0=1'h0;
wire	[1:0]	mux_u104_u0;
wire		or_u372_u0;
wire		mux_u105_u0;
wire		or_u373_u0;
wire	[31:0]	mux_u106_u0;
wire		or_u374_u0;
wire		or_u375_u0;
wire	[31:0]	mux_u107_u0;
wire	[1:0]	mux_u108_u0;
wire		or_u376_u0;
reg		reg_65426ec1_result_delayed_u0=1'h0;
assign and_u1341_u0=or_u371_u0&or_u371_u0;
assign equals_a_signed=port_2b235147_;
assign equals_b_signed=32'h40000;
assign equals=equals_a_signed==equals_b_signed;
assign equals_u74_a_signed=port_2b235147_;
assign equals_u74_b_signed=32'h40000;
assign equals_u74=equals_u74_a_signed==equals_u74_b_signed;
assign equals_u75_a_signed=port_5b5cde36_;
assign equals_u75_b_signed=32'h2;
assign equals_u75=equals_u75_a_signed==equals_u75_b_signed;
assign equals_u76_a_signed={30'b0, syncEnable_u89_u0[1:0]};
assign equals_u76_b_signed=32'h0;
assign equals_u76=equals_u76_a_signed==equals_u76_b_signed;
assign and_u1342_u0=block_GO_delayed_u1_u0&equals_u76;
assign and_u1343_u0=block_GO_delayed_u1_u0&not_u255_u0;
assign not_u255_u0=~equals_u76;
assign and_u1344_u0=and_u1349_u0&syncEnable_u83_u0;
assign not_u256_u0=~syncEnable_u83_u0;
assign and_u1345_u0=and_u1349_u0&not_u256_u0;
assign simplePinWrite=and_u1347_u0&{1{and_u1347_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_55828783_u0<=1'h0;
else reg_55828783_u0<=and_u1346_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_39bf2b99_u0<=1'h0;
else reg_39bf2b99_u0<=and_u1347_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_39bf2b99_result_delayed_u0<=1'h0;
else reg_39bf2b99_result_delayed_u0<=reg_39bf2b99_u0;
end
assign and_u1346_u0=and_u1345_u0&and_u1349_u0;
assign or_u349_u0=reg_55828783_u0|reg_39bf2b99_result_delayed_result_delayed_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_39bf2b99_result_delayed_result_delayed_u0<=1'h0;
else reg_39bf2b99_result_delayed_result_delayed_u0<=reg_39bf2b99_result_delayed_u0;
end
assign and_u1347_u0=and_u1344_u0&and_u1349_u0;
assign mux_u88=(and_u1347_u0)?2'h1:2'h3;
assign or_u350_u0=and_u1347_u0|and_u1346_u0;
assign or_u351_u0=and_delayed_u71|or_u349_u0;
assign and_u1348_u0=and_u1343_u0&block_GO_delayed_u1_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u71<=1'h0;
else and_delayed_u71<=and_u1348_u0;
end
assign and_u1349_u0=and_u1342_u0&block_GO_delayed_u1_u0;
assign equals_u77_a_signed={30'b0, syncEnable_u89_u0[1:0]};
assign equals_u77_b_signed=32'h1;
assign equals_u77=equals_u77_a_signed==equals_u77_b_signed;
assign not_u257_u0=~equals_u77;
assign and_u1350_u0=block_GO_delayed_u1_u0&equals_u77;
assign and_u1351_u0=block_GO_delayed_u1_u0&not_u257_u0;
assign and_u1352_u0=and_u1368_u0&syncEnable_u88_u0;
assign and_u1353_u0=and_u1368_u0&not_u258_u0;
assign not_u258_u0=~syncEnable_u88_u0;
assign andOp=port_01ffd1e5_&port_2d451d49_;
assign not_u259_u0=~andOp;
assign and_u1354_u0=and_u1366_u0&not_u259_u0;
assign and_u1355_u0=and_u1366_u0&andOp;
assign simplePinWrite_u223=and_u1356_u0&{1{and_u1356_u0}};
assign or_u352_u0=reg_49e39485_u0|and_delayed_u73_u0;
assign and_u1356_u0=and_u1355_u0&and_u1366_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_49e39485_u0<=1'h0;
else reg_49e39485_u0<=and_delayed_u72_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u72_u0<=1'h0;
else and_delayed_u72_u0<=and_u1356_u0;
end
assign and_u1357_u0=and_u1354_u0&and_u1366_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u73_u0<=1'h0;
else and_delayed_u73_u0<=and_u1357_u0;
end
assign and_u1358_u0=and_u1367_u0&not_u260_u0;
assign not_u260_u0=~syncEnable_u85_u0;
assign and_u1359_u0=and_u1367_u0&syncEnable_u85_u0;
assign and_u1360_u0=and_u1364_u0&port_2d451d49_;
assign not_u261_u0=~port_2d451d49_;
assign and_u1361_u0=and_u1364_u0&not_u261_u0;
assign simplePinWrite_u224=and_u1362_u0&{1{and_u1362_u0}};
assign or_u353_u0=reg_64307160_u0|reg_7a1ee0d6_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a1ee0d6_u0<=1'h0;
else reg_7a1ee0d6_u0<=reg_7bb2e7de_u0;
end
assign and_u1362_u0=and_u1360_u0&and_u1364_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7bb2e7de_u0<=1'h0;
else reg_7bb2e7de_u0<=and_delayed_u74_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_64307160_u0<=1'h0;
else reg_64307160_u0<=and_u1363_u0;
end
assign and_u1363_u0=and_u1361_u0&and_u1364_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u74_u0<=1'h0;
else and_delayed_u74_u0<=and_u1362_u0;
end
assign and_u1364_u0=and_u1359_u0&and_u1367_u0;
assign or_u354_u0=and_delayed_u75_u0|or_u353_u0;
assign and_u1365_u0=and_u1358_u0&and_u1367_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u75_u0<=1'h0;
else and_delayed_u75_u0<=and_u1365_u0;
end
assign mux_u89_u0=(and_u1362_u0)?2'h2:2'h3;
assign or_u355_u0=and_u1362_u0|and_u1365_u0;
assign or_u356_u0=or_u352_u0|or_u354_u0;
assign mux_u90_u0=(and_u1356_u0)?2'h0:{1'b1, mux_u89_u0[0]};
assign or_u357_u0=and_u1356_u0|or_u355_u0;
assign and_u1366_u0=and_u1352_u0&and_u1368_u0;
assign and_u1367_u0=and_u1353_u0&and_u1368_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00382bbc_u0<=1'h0;
else reg_00382bbc_u0<=and_u1369_u0;
end
assign and_u1368_u0=and_u1350_u0&block_GO_delayed_u1_u0;
assign or_u358_u0=or_u356_u0|reg_00382bbc_u0;
assign and_u1369_u0=and_u1351_u0&block_GO_delayed_u1_u0;
assign equals_u78_a_signed={30'b0, syncEnable_u89_u0[1:0]};
assign equals_u78_b_signed=32'h2;
assign equals_u78=equals_u78_a_signed==equals_u78_b_signed;
assign and_u1370_u0=block_GO_delayed_u1_u0&equals_u78;
assign and_u1371_u0=block_GO_delayed_u1_u0&not_u262_u0;
assign not_u262_u0=~equals_u78;
assign and_u1372_u0=and_u1389_u0&not_u263_u0;
assign not_u263_u0=~syncEnable_u90_u0;
assign and_u1373_u0=and_u1389_u0&syncEnable_u90_u0;
assign andOp_u108=port_01ffd1e5_&port_2d451d49_;
assign and_u1374_u0=and_u1387_u0&andOp_u108;
assign not_u264_u0=~andOp_u108;
assign and_u1375_u0=and_u1387_u0&not_u264_u0;
assign simplePinWrite_u225=and_u1376_u0&{1{and_u1376_u0}};
assign and_u1376_u0=and_u1374_u0&and_u1387_u0;
assign and_u1377_u0=and_u1375_u0&and_u1387_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_04ddc90f_u0<=1'h0;
else reg_04ddc90f_u0<=and_delayed_u77_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u76_u0<=1'h0;
else and_delayed_u76_u0<=and_u1377_u0;
end
assign or_u359_u0=reg_04ddc90f_u0|and_delayed_u76_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u77_u0<=1'h0;
else and_delayed_u77_u0<=and_u1376_u0;
end
assign not_u265_u0=~syncEnable_u92_u0;
assign and_u1378_u0=and_u1386_u0&syncEnable_u92_u0;
assign and_u1379_u0=and_u1386_u0&not_u265_u0;
assign and_u1380_u0=and_u1385_u0&port_01ffd1e5_;
assign not_u266_u0=~port_01ffd1e5_;
assign and_u1381_u0=and_u1385_u0&not_u266_u0;
assign simplePinWrite_u226=and_u1383_u0&{1{and_u1383_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5ed9e738_u0<=1'h0;
else reg_5ed9e738_u0<=and_u1383_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_679f5f5d_u0<=1'h0;
else reg_679f5f5d_u0<=reg_5ed9e738_result_delayed_u0;
end
assign or_u360_u0=reg_679f5f5d_u0|and_delayed_u78_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5ed9e738_result_delayed_u0<=1'h0;
else reg_5ed9e738_result_delayed_u0<=reg_5ed9e738_u0;
end
assign and_u1382_u0=and_u1381_u0&and_u1385_u0;
assign and_u1383_u0=and_u1380_u0&and_u1385_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u78_u0<=1'h0;
else and_delayed_u78_u0<=and_u1382_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5cab12fe_u0<=1'h0;
else reg_5cab12fe_u0<=and_u1384_u0;
end
assign and_u1384_u0=and_u1379_u0&and_u1386_u0;
assign or_u361_u0=reg_5cab12fe_u0|or_u360_u0;
assign mux_u91_u0=(and_u1383_u0)?2'h1:2'h3;
assign or_u362_u0=and_u1383_u0|and_u1384_u0;
assign and_u1385_u0=and_u1378_u0&and_u1386_u0;
assign and_u1386_u0=and_u1372_u0&and_u1389_u0;
assign and_u1387_u0=and_u1373_u0&and_u1389_u0;
assign or_u363_u0=or_u359_u0|or_u361_u0;
assign or_u364_u0=and_u1376_u0|or_u362_u0;
assign mux_u92_u0=(and_u1376_u0)?2'h0:{mux_u91_u0[1], 1'b1};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_29f791b4_u0<=1'h0;
else reg_29f791b4_u0<=and_u1388_u0;
end
assign and_u1388_u0=and_u1371_u0&block_GO_delayed_u1_u0;
assign or_u365_u0=or_u363_u0|reg_29f791b4_u0;
assign and_u1389_u0=and_u1370_u0&block_GO_delayed_u1_u0;
assign equals_u79_a_signed={30'b0, syncEnable_u89_u0[1:0]};
assign equals_u79_b_signed=32'h3;
assign equals_u79=equals_u79_a_signed==equals_u79_b_signed;
assign and_u1390_u0=block_GO_delayed_u1_u0&not_u267_u0;
assign and_u1391_u0=block_GO_delayed_u1_u0&equals_u79;
assign not_u267_u0=~equals_u79;
assign lessThan_a_signed=syncEnable_u87_u0;
assign lessThan_b_signed=syncEnable_u91_u0;
assign lessThan=lessThan_a_signed<lessThan_b_signed;
assign not_u268_u0=~lessThan;
assign and_u1392_u0=and_u1401_u0&not_u268_u0;
assign and_u1393_u0=and_u1401_u0&lessThan;
assign and_u1394_u0=and_u1400_u0&syncEnable_u84_u0;
assign not_u269_u0=~syncEnable_u84_u0;
assign and_u1395_u0=and_u1400_u0&not_u269_u0;
assign simplePinWrite_u227=and_u1397_u0&{1{and_u1397_u0}};
assign add=syncEnable_u87_u0+32'h0;
always @(posedge CLK or posedge and_u1397_u0 or posedge or_u366_u0)
begin
if (or_u366_u0)
reg_22328357_u0<=1'h0;
else if (and_u1397_u0)
reg_22328357_u0<=1'h1;
else reg_22328357_u0<=reg_22328357_u0;
end
assign or_u366_u0=and_u1396_u0|RESET;
assign and_u1396_u0=reg_22328357_u0&port_30bf0bb1_;
assign add_u33=syncEnable_u87_u0+32'h1;
always @(posedge CLK)
begin
if (and_u1397_u0)
syncEnable_u76<=port_7dc7ca1e_;
end
assign and_u1397_u0=and_u1394_u0&and_u1400_u0;
assign mux_u93_u0=(and_delayed_u79_u0)?syncEnable_u76:syncEnable_u77_u0;
assign and_u1398_u0=and_u1395_u0&and_u1400_u0;
always @(posedge CLK)
begin
if (and_u1400_u0)
syncEnable_u77_u0<=syncEnable_u93_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u79_u0<=1'h0;
else and_delayed_u79_u0<=and_u1397_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u80_u0<=1'h0;
else and_delayed_u80_u0<=and_u1398_u0;
end
always @(posedge CLK)
begin
if (and_u1399_u0)
syncEnable_u78_u0<={1'b0, port_18e00d02_};
end
always @(posedge CLK)
begin
if (and_u1401_u0)
syncEnable_u79_u0<=syncEnable_u93_u0;
end
assign and_u1399_u0=and_u1392_u0&and_u1401_u0;
assign mux_u94_u0=(and_delayed_u81_u0)?mux_u93_u0:syncEnable_u79_u0;
always @(posedge CLK)
begin
if (and_u1401_u0)
syncEnable_u80_u0<=syncEnable_u86_u0;
end
assign and_u1400_u0=and_u1393_u0&and_u1401_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u81_u0<=1'h0;
else and_delayed_u81_u0<=and_u1400_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u82_u0<=1'h0;
else and_delayed_u82_u0<=and_u1399_u0;
end
assign mux_u95_u0=(and_delayed_u81_u0)?syncEnable_u80_u0:{30'b0, syncEnable_u78_u0[1:0]};
assign mux_u96_u0=(and_delayed_u83_u0)?mux_u94_u0:syncEnable_u81_u0;
assign mux_u97_u0=(and_delayed_u83_u0)?mux_u95_u0:syncEnable_u82_u0;
assign and_u1401_u0=and_u1391_u0&block_GO_delayed_u1_u0;
assign and_u1402_u0=and_u1390_u0&block_GO_delayed_u1_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u83_u0<=1'h0;
else and_delayed_u83_u0<=and_u1401_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u84_u0<=1'h0;
else and_delayed_u84_u0<=and_u1402_u0;
end
always @(posedge CLK)
begin
if (block_GO_delayed_u1_u0)
syncEnable_u81_u0<=syncEnable_u93_u0;
end
always @(posedge CLK)
begin
if (block_GO_delayed_u1_u0)
syncEnable_u82_u0<=syncEnable_u86_u0;
end
assign latch_1f7403f6_out=(block_GO_delayed_u0)?mux_u97_u0:latch_1f7403f6_reg;
always @(posedge CLK)
begin
if (block_GO_delayed_u0)
latch_1f7403f6_reg<=mux_u97_u0;
end
assign or_u367_u0=and_u1346_u0|and_u1399_u0;
assign mux_u98_u0=(and_u1346_u0)?32'h0:32'hfffffffd;
assign or_u368_u0=and_u1346_u0|and_u1365_u0|and_u1384_u0;
assign mux_u99_u0=({2{and_u1346_u0}}&2'h0)|({2{and_u1365_u0}}&2'h1)|({2{and_u1384_u0}}&2'h2);
assign mux_u100_u0=({2{or_u350_u0}}&{mux_u88[1], 1'b1})|({2{or_u357_u0}}&mux_u90_u0)|({2{or_u364_u0}}&mux_u92_u0)|({2{and_u1399_u0}}&port_18e00d02_);
assign or_u369_u0=or_u350_u0|or_u357_u0|or_u364_u0|and_u1399_u0;
assign or_u370_u0=and_u1347_u0|and_u1397_u0;
assign mux_u101_u0=(and_u1347_u0)?32'h0:add_u33;
always @(posedge CLK)
begin
if (bus_3c51dea1_)
scoreboard_428a1a5c_reg1<=1'h0;
else if (or_u365_u0)
scoreboard_428a1a5c_reg1<=1'h1;
else scoreboard_428a1a5c_reg1<=scoreboard_428a1a5c_reg1;
end
assign scoreboard_428a1a5c_resOr0=or_u351_u0|scoreboard_428a1a5c_reg0;
assign scoreboard_428a1a5c_and=scoreboard_428a1a5c_resOr0&scoreboard_428a1a5c_resOr1&scoreboard_428a1a5c_resOr2;
assign scoreboard_428a1a5c_resOr1=or_u365_u0|scoreboard_428a1a5c_reg1;
assign bus_3c51dea1_=scoreboard_428a1a5c_and|RESET;
always @(posedge CLK)
begin
if (bus_3c51dea1_)
scoreboard_428a1a5c_reg0<=1'h0;
else if (or_u351_u0)
scoreboard_428a1a5c_reg0<=1'h1;
else scoreboard_428a1a5c_reg0<=scoreboard_428a1a5c_reg0;
end
always @(posedge CLK)
begin
if (bus_3c51dea1_)
scoreboard_428a1a5c_reg2<=1'h0;
else if (or_u358_u0)
scoreboard_428a1a5c_reg2<=1'h1;
else scoreboard_428a1a5c_reg2<=scoreboard_428a1a5c_reg2;
end
assign scoreboard_428a1a5c_resOr2=or_u358_u0|scoreboard_428a1a5c_reg2;
always @(posedge CLK)
begin
if (block_GO_delayed_u0)
latch_7da74311_reg<=mux_u96_u0;
end
assign latch_7da74311_out=(block_GO_delayed_u0)?mux_u96_u0:latch_7da74311_reg;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
block_GO_delayed_u0<=1'h0;
else block_GO_delayed_u0<=block_GO_delayed_u1_u0;
end
always @(posedge CLK)
begin
if (and_u1341_u0)
syncEnable_u83_u0<=equals_u75;
end
always @(posedge CLK)
begin
if (and_u1341_u0)
syncEnable_u84_u0<=port_2cc0cc2a_;
end
always @(posedge CLK)
begin
if (and_u1341_u0)
syncEnable_u85_u0<=port_2cc0cc2a_;
end
always @(posedge CLK)
begin
if (and_u1341_u0)
syncEnable_u86_u0<=mux_u103_u0;
end
always @(posedge CLK)
begin
if (and_u1341_u0)
syncEnable_u87_u0<=port_5b5cde36_;
end
always @(posedge CLK)
begin
if (and_u1341_u0)
syncEnable_u88_u0<=equals;
end
always @(posedge CLK)
begin
if (and_u1341_u0)
syncEnable_u89_u0<={1'b0, port_7b9868d2_};
end
always @(posedge CLK)
begin
if (and_u1341_u0)
syncEnable_u90_u0<=equals_u74;
end
always @(posedge CLK)
begin
if (and_u1341_u0)
syncEnable_u91_u0<=port_7a3e2d5e_;
end
always @(posedge CLK)
begin
if (and_u1341_u0)
syncEnable_u92_u0<=port_2cc0cc2a_;
end
always @(posedge CLK)
begin
if (and_u1341_u0)
syncEnable_u93_u0<=mux_u102_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
block_GO_delayed_u1_u0<=1'h0;
else block_GO_delayed_u1_u0<=and_u1341_u0;
end
assign mux_u102_u0=(loopControl_u0)?fbReg_In1Portvalue_u0:16'h0;
always @(posedge CLK)
begin
if (scoreboard_428a1a5c_and)
fbReg_temp_fsmOldState_image1_iunzip_0_u0<=latch_1f7403f6_out;
end
always @(posedge CLK)
begin
if (scoreboard_428a1a5c_and)
fbReg_In1Portvalue_u0<=latch_7da74311_out;
end
always @(posedge CLK)
begin
if (reg_65426ec1_result_delayed_u0)
syncEnable_u94_u0<=RESET;
end
always @(posedge CLK or posedge syncEnable_u94_u0)
begin
if (syncEnable_u94_u0)
loopControl_u0<=1'h0;
else loopControl_u0<=scoreboard_428a1a5c_and;
end
assign or_u371_u0=loopControl_u0|reg_65426ec1_result_delayed_u0;
assign mux_u103_u0=(loopControl_u0)?fbReg_temp_fsmOldState_image1_iunzip_0_u0:32'h0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_65426ec1_u0<=1'h0;
else reg_65426ec1_u0<=GO;
end
assign mux_u104_u0=(GO)?2'h0:mux_u99_u0;
assign or_u372_u0=GO|or_u368_u0;
assign mux_u105_u0=(GO)?1'h0:1'h1;
assign or_u373_u0=GO|and_u1346_u0;
assign mux_u106_u0=(GO)?32'h0:mux_u101_u0;
assign or_u374_u0=GO|or_u370_u0;
assign or_u375_u0=GO|or_u367_u0;
assign mux_u107_u0=(GO)?32'hfffffffd:{mux_u98_u0[31:2], 1'b0, mux_u98_u0[0]};
assign mux_u108_u0=(GO)?2'h0:mux_u100_u0;
assign or_u376_u0=GO|or_u369_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_65426ec1_result_delayed_u0<=1'h0;
else reg_65426ec1_result_delayed_u0<=reg_65426ec1_u0;
end
assign RESULT=or_u372_u0;
assign RESULT_u787=mux_u104_u0;
assign RESULT_u788=or_u376_u0;
assign RESULT_u789=mux_u108_u0;
assign RESULT_u790=or_u374_u0;
assign RESULT_u791=mux_u106_u0;
assign RESULT_u792=or_u375_u0;
assign RESULT_u793={mux_u107_u0[31:2], 1'b0, mux_u107_u0[0]};
assign RESULT_u794=or_u373_u0;
assign RESULT_u795=mux_u105_u0;
assign RESULT_u796=and_u1397_u0;
assign RESULT_u797=add;
assign RESULT_u798=port_7dc7ca1e_;
assign RESULT_u799=3'h1;
assign RESULT_u800=simplePinWrite;
assign RESULT_u801=simplePinWrite_u224;
assign RESULT_u802=simplePinWrite_u226;
assign RESULT_u803=simplePinWrite_u225;
assign RESULT_u804=simplePinWrite_u227;
assign RESULT_u805=simplePinWrite_u223;
assign DONE=1'h0;
endmodule



module image1_iunzip_simplememoryreferee_3f8b2b7e_(bus_4fdc6d9e_, bus_16db627b_, bus_5c6b1ef6_, bus_7e5a1f5a_, bus_220ac51f_, bus_77abea3c_, bus_55f9978e_, bus_192ef9bb_, bus_26fb90a8_, bus_5ac8d702_, bus_5fd8a7cf_, bus_73bd858d_, bus_592fb24a_, bus_68afb47e_, bus_1604219b_, bus_7a726660_, bus_4ba2e658_, bus_394326ad_, bus_4399e227_);
input		bus_4fdc6d9e_;
input		bus_16db627b_;
input		bus_5c6b1ef6_;
input	[15:0]	bus_7e5a1f5a_;
input		bus_220ac51f_;
input	[31:0]	bus_77abea3c_;
input	[2:0]	bus_55f9978e_;
input		bus_192ef9bb_;
input	[15:0]	bus_26fb90a8_;
input	[31:0]	bus_5ac8d702_;
input	[2:0]	bus_5fd8a7cf_;
output	[15:0]	bus_73bd858d_;
output	[31:0]	bus_592fb24a_;
output		bus_68afb47e_;
output		bus_1604219b_;
output	[2:0]	bus_7a726660_;
output	[15:0]	bus_4ba2e658_;
output		bus_394326ad_;
output		bus_4399e227_;
reg		done_qual_u46_u0=1'h0;
wire		or_6aa3cfa4_u0;
wire		or_7cc2a2ea_u0;
wire		or_596c9963_u0;
wire		not_3181d6ce_u0;
wire		and_11031633_u0;
wire	[31:0]	mux_5f778cc6_u0;
wire	[15:0]	mux_1a840f9e_u0;
wire		and_47c44019_u0;
wire		not_4252c80c_u0;
reg		done_qual_u47_u0=1'h0;
always @(posedge bus_4fdc6d9e_)
begin
if (bus_16db627b_)
done_qual_u46_u0<=1'h0;
else done_qual_u46_u0<=bus_220ac51f_;
end
assign or_6aa3cfa4_u0=bus_192ef9bb_|done_qual_u47_u0;
assign or_7cc2a2ea_u0=bus_220ac51f_|done_qual_u46_u0;
assign bus_73bd858d_=mux_1a840f9e_u0;
assign bus_592fb24a_=mux_5f778cc6_u0;
assign bus_68afb47e_=bus_192ef9bb_;
assign bus_1604219b_=or_596c9963_u0;
assign bus_7a726660_=3'h1;
assign bus_4ba2e658_=bus_7e5a1f5a_;
assign bus_394326ad_=and_11031633_u0;
assign bus_4399e227_=and_47c44019_u0;
assign or_596c9963_u0=bus_220ac51f_|bus_192ef9bb_;
assign not_3181d6ce_u0=~bus_5c6b1ef6_;
assign and_11031633_u0=or_7cc2a2ea_u0&bus_5c6b1ef6_;
assign mux_5f778cc6_u0=(bus_220ac51f_)?32'h0:bus_5ac8d702_;
assign mux_1a840f9e_u0=({16{bus_192ef9bb_}}&bus_26fb90a8_);
assign and_47c44019_u0=or_6aa3cfa4_u0&bus_5c6b1ef6_;
assign not_4252c80c_u0=~bus_5c6b1ef6_;
always @(posedge bus_4fdc6d9e_)
begin
if (bus_16db627b_)
done_qual_u47_u0<=1'h0;
else done_qual_u47_u0<=bus_192ef9bb_;
end
endmodule



module image1_iunzip_globalreset_physical_0787df71_(bus_137e2708_, bus_19659027_, bus_5857bbf3_);
input		bus_137e2708_;
input		bus_19659027_;
output		bus_5857bbf3_;
wire		and_167aac1b_u0;
reg		final_u18=1'h1;
reg		glitch_u18=1'h0;
wire		or_298f8509_u0;
reg		sample_u18=1'h0;
wire		not_1ef482b8_u0;
reg		cross_u18=1'h0;
assign and_167aac1b_u0=cross_u18&glitch_u18;
always @(posedge bus_137e2708_)
begin
final_u18<=not_1ef482b8_u0;
end
assign bus_5857bbf3_=or_298f8509_u0;
always @(posedge bus_137e2708_)
begin
glitch_u18<=cross_u18;
end
assign or_298f8509_u0=bus_19659027_|final_u18;
always @(posedge bus_137e2708_)
begin
sample_u18<=1'h1;
end
assign not_1ef482b8_u0=~and_167aac1b_u0;
always @(posedge bus_137e2708_)
begin
cross_u18<=sample_u18;
end
endmodule



module image1_iunzip_forge_memory_3x16_7(CLK, ENA, WEA, DINA, ENB, ADDRA, ADDRB, DOUTA, DOUTB, DONEA, DONEB);
input		CLK;
input		ENA;
input		WEA;
input	[15:0]	DINA;
input		ENB;
input	[31:0]	ADDRA;
input	[31:0]	ADDRB;
output	[15:0]	DOUTA;
output	[15:0]	DOUTB;
output		DONEA;
output		DONEB;
wire		wea_0;
wire	[15:0]	pre_douta_0;
wire	[15:0]	pre_doutb_0;
reg		wea_done;
reg		rea_done;
reg	[15:0]	mux_outa;
reg	[15:0]	mux_outb;
assign wea_0=WEA;
always @(posedge CLK)
begin
wea_done<=WEA;
end
assign DONEA=rea_done|wea_done;
always @(posedge CLK)
begin
end
assign DONEB=ENB;
always @(pre_douta_0)
begin
mux_outa<=pre_douta_0;
end
assign DOUTA=mux_outa;
always @(pre_doutb_0)
begin
mux_outb<=pre_doutb_0;
end
assign DOUTB=mux_outb;
// Memory array element: COL: 0, ROW: 0
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_16(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[0]), .SPO(pre_douta_0[0]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[0]));
// Memory array element: COL: 0, ROW: 1
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_17(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[1]), .SPO(pre_douta_0[1]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[1]));
// Memory array element: COL: 0, ROW: 2
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_18(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[2]), .SPO(pre_douta_0[2]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[2]));
// Memory array element: COL: 0, ROW: 3
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_19(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[3]), .SPO(pre_douta_0[3]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[3]));
// Memory array element: COL: 0, ROW: 4
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_20(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[4]), .SPO(pre_douta_0[4]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[4]));
// Memory array element: COL: 0, ROW: 5
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_21(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[5]), .SPO(pre_douta_0[5]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[5]));
// Memory array element: COL: 0, ROW: 6
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_22(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[6]), .SPO(pre_douta_0[6]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[6]));
// Memory array element: COL: 0, ROW: 7
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_23(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[7]), .SPO(pre_douta_0[7]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[7]));
// Memory array element: COL: 0, ROW: 8
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_24(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[8]), .SPO(pre_douta_0[8]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[8]));
// Memory array element: COL: 0, ROW: 9
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_25(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[9]), .SPO(pre_douta_0[9]), .DPRA0(ADDRB[0]), 
  .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[9]));
// Memory array element: COL: 0, ROW: 10
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_26(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[10]), .SPO(pre_douta_0[10]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[10]));
// Memory array element: COL: 0, ROW: 11
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_27(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[11]), .SPO(pre_douta_0[11]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[11]));
// Memory array element: COL: 0, ROW: 12
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_28(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[12]), .SPO(pre_douta_0[12]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[12]));
// Memory array element: COL: 0, ROW: 13
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_29(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[13]), .SPO(pre_douta_0[13]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[13]));
// Memory array element: COL: 0, ROW: 14
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_30(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[14]), .SPO(pre_douta_0[14]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[14]));
// Memory array element: COL: 0, ROW: 15
//  Initialization of Dual Port LUT ram now done through explicit
// parameter setting.
RAM16X1D#(.INIT(16'h0000))RAM16X1D_instance_31(.WCLK(CLK), .WE(wea_0), .A0(ADDRA[0]), 
  .A1(ADDRA[1]), .A2(ADDRA[2]), .A3(ADDRA[3]), .D(DINA[15]), .SPO(pre_douta_0[15]), 
  .DPRA0(ADDRB[0]), .DPRA1(ADDRB[1]), .DPRA2(ADDRB[2]), .DPRA3(ADDRB[3]), .DPO(pre_doutb_0[15]));
endmodule



module image1_iunzip_structuralmemory_224e8538_(CLK_u3, bus_44b4fa91_, bus_0f1d20b4_, bus_625040d8_, bus_38cab4e5_, bus_1f7bdd2e_, bus_4944043d_, bus_2448127a_, bus_016e260c_, bus_25f12fe5_, bus_6d3e7bde_, bus_6204046f_, bus_0c649092_, bus_4cc7a537_);
input		CLK_u3;
input		bus_44b4fa91_;
input	[31:0]	bus_0f1d20b4_;
input	[2:0]	bus_625040d8_;
input		bus_38cab4e5_;
input		bus_1f7bdd2e_;
input	[15:0]	bus_4944043d_;
input	[31:0]	bus_2448127a_;
input	[2:0]	bus_016e260c_;
input		bus_25f12fe5_;
output	[15:0]	bus_6d3e7bde_;
output		bus_6204046f_;
output	[15:0]	bus_0c649092_;
output		bus_4cc7a537_;
wire		not_43a4e7ce_u0;
wire		or_1ed5ab5a_u0;
wire		and_523a7468_u0;
wire		or_4a23b6b4_u0;
wire	[15:0]	bus_0b1d7167_;
wire	[15:0]	bus_289877c2_;
reg		logicalMem_6aebccf8_we_delay0_u0=1'h0;
assign not_43a4e7ce_u0=~bus_1f7bdd2e_;
assign or_1ed5ab5a_u0=and_523a7468_u0|logicalMem_6aebccf8_we_delay0_u0;
assign and_523a7468_u0=bus_38cab4e5_&not_43a4e7ce_u0;
assign or_4a23b6b4_u0=bus_38cab4e5_|bus_1f7bdd2e_;
image1_iunzip_forge_memory_3x16_7 image1_iunzip_forge_memory_3x16_7_instance0(.CLK(CLK_u3), 
  .ENA(or_4a23b6b4_u0), .WEA(bus_1f7bdd2e_), .DINA(bus_4944043d_), .ADDRA(bus_0f1d20b4_), 
  .DOUTA(bus_289877c2_), .DONEA(), .ENB(bus_25f12fe5_), .ADDRB(bus_2448127a_), .DOUTB(bus_0b1d7167_), 
  .DONEB());
assign bus_6d3e7bde_=bus_289877c2_;
assign bus_6204046f_=or_1ed5ab5a_u0;
assign bus_0c649092_=bus_0b1d7167_;
assign bus_4cc7a537_=bus_25f12fe5_;
always @(posedge CLK_u3 or posedge bus_44b4fa91_)
begin
if (bus_44b4fa91_)
logicalMem_6aebccf8_we_delay0_u0<=1'h0;
else logicalMem_6aebccf8_we_delay0_u0<=bus_1f7bdd2e_;
end
endmodule



module image1_iunzip_streamEndFun2(CLK, RESET, GO, port_63ac392a_, port_4739a893_, port_2068be2c_, port_1e8c51ba_, port_177ce6b0_, RESULT, RESULT_u806, RESULT_u807, RESULT_u808, RESULT_u809, RESULT_u810, RESULT_u811, RESULT_u812, RESULT_u813, RESULT_u814, RESULT_u815, RESULT_u816, RESULT_u817, RESULT_u818, DONE);
input		CLK;
input		RESET;
input		GO;
input		port_63ac392a_;
input		port_4739a893_;
input	[15:0]	port_2068be2c_;
input		port_1e8c51ba_;
input	[15:0]	port_177ce6b0_;
output		RESULT;
output		RESULT_u806;
output		RESULT_u807;
output	[31:0]	RESULT_u808;
output	[2:0]	RESULT_u809;
output		RESULT_u810;
output	[31:0]	RESULT_u811;
output	[2:0]	RESULT_u812;
output	[15:0]	RESULT_u813;
output	[15:0]	RESULT_u814;
output		RESULT_u815;
output		RESULT_u816;
output	[15:0]	RESULT_u817;
output	[15:0]	RESULT_u818;
output		DONE;
wire	[31:0]	add;
wire		and_u1403_u0;
wire	[8:0]	subtract;
wire signed	[8:0]	greaterThanEqualTo_b_signed;
wire signed	[8:0]	greaterThanEqualTo_a_signed;
wire		greaterThanEqualTo;
wire		and_u1404_u0;
wire		not_u270_u0;
wire		and_u1405_u0;
wire	[8:0]	subtract_u5;
wire		and_u1406_u0;
wire	[8:0]	mux_u109;
wire		and_u1407_u0;
wire	[31:0]	add_u34;
wire		and_u1408_u0;
wire		and_u1410_u0;
wire	[16:0]	add_u35;
wire	[15:0]	add_u36;
wire	[15:0]	simplePinWrite;
wire	[15:0]	simplePinWrite_u228;
wire		simplePinWrite_u229;
wire	[15:0]	simplePinWrite_u230;
wire		simplePinWrite_u231;
wire	[15:0]	simplePinWrite_u232;
reg	[31:0]	syncEnable_u95=32'h0;
reg	[15:0]	syncEnable_u96_u0=16'h0;
wire		or_u377_u0;
wire	[31:0]	mux_u110_u0;
reg		reg_4fbb82fa_u0=1'h0;
reg	[31:0]	syncEnable_u97_u0=32'h0;
reg	[15:0]	syncEnable_u98_u0=16'h0;
reg		reg_4fbb82fa_result_delayed_u0=1'h0;
assign add={31'b0, port_63ac392a_}+32'h0;
assign and_u1403_u0=reg_4fbb82fa_u0&port_1e8c51ba_;
assign subtract={8'b0, port_63ac392a_}-9'h1;
assign greaterThanEqualTo_a_signed={subtract[2], subtract[2], subtract[2], subtract[2], subtract[2], subtract[2], subtract[2:0]};
assign greaterThanEqualTo_b_signed=9'h0;
assign greaterThanEqualTo=greaterThanEqualTo_a_signed>=greaterThanEqualTo_b_signed;
assign and_u1404_u0=GO&greaterThanEqualTo;
assign not_u270_u0=~greaterThanEqualTo;
assign and_u1405_u0=GO&not_u270_u0;
assign subtract_u5={8'b0, port_63ac392a_}-9'h1;
assign and_u1406_u0=and_u1404_u0&GO;
assign mux_u109=(and_u1406_u0)?{subtract_u5[2], subtract_u5[2], subtract_u5[2], subtract_u5[2], subtract_u5[2], subtract_u5[2], subtract_u5[2:0]}:9'h2;
assign and_u1407_u0=and_u1405_u0&GO;
assign add_u34={mux_u109[2], mux_u109[2], mux_u109[2], mux_u109[2], mux_u109[2], mux_u109[2], mux_u109[2], mux_u109[2], mux_u109[2], mux_u109[2], mux_u109[2], mux_u109[2], mux_u109[2], mux_u109[2], mux_u109[2], mux_u109[2], mux_u109[2], mux_u109[2], mux_u109[2], mux_u109[2], mux_u109[2], mux_u109[2], mux_u109[2], mux_u109[2], mux_u109[2], mux_u109[2], mux_u109[2], mux_u109[2], mux_u109[2], mux_u109[2:0]}+32'h0;
assign and_u1408_u0=reg_4fbb82fa_u0&port_4739a893_;
assign and_u1410_u0=reg_4fbb82fa_result_delayed_u0&port_1e8c51ba_;
assign add_u35={syncEnable_u96_u0[15], syncEnable_u96_u0}+{port_177ce6b0_[15], port_177ce6b0_};
assign add_u36=syncEnable_u98_u0+{add_u35[16], add_u35[16:2]};
assign simplePinWrite=add_u36&{16{reg_4fbb82fa_result_delayed_u0}};
assign simplePinWrite_u228=16'h1&{16{1'h1}};
assign simplePinWrite_u229=reg_4fbb82fa_result_delayed_u0&{1{reg_4fbb82fa_result_delayed_u0}};
assign simplePinWrite_u230=16'h1&{16{1'h1}};
assign simplePinWrite_u231=reg_4fbb82fa_result_delayed_u0&{1{reg_4fbb82fa_result_delayed_u0}};
assign simplePinWrite_u232=add_u36&{16{reg_4fbb82fa_result_delayed_u0}};
always @(posedge CLK)
begin
if (GO)
syncEnable_u95<={add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2], add[2:0]};
end
always @(posedge CLK)
begin
if (reg_4fbb82fa_u0)
syncEnable_u96_u0<=port_2068be2c_;
end
assign or_u377_u0=reg_4fbb82fa_u0|reg_4fbb82fa_result_delayed_u0;
assign mux_u110_u0=(reg_4fbb82fa_u0)?syncEnable_u95:32'h0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4fbb82fa_u0<=1'h0;
else reg_4fbb82fa_u0<=GO;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u97_u0<=add_u34;
end
always @(posedge CLK)
begin
if (reg_4fbb82fa_u0)
syncEnable_u98_u0<=port_177ce6b0_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4fbb82fa_result_delayed_u0<=1'h0;
else reg_4fbb82fa_result_delayed_u0<=reg_4fbb82fa_u0;
end
assign RESULT=GO;
assign RESULT_u806=1'h0;
assign RESULT_u807=reg_4fbb82fa_u0;
assign RESULT_u808=syncEnable_u97_u0;
assign RESULT_u809=3'h1;
assign RESULT_u810=or_u377_u0;
assign RESULT_u811=mux_u110_u0;
assign RESULT_u812=3'h1;
assign RESULT_u813=simplePinWrite_u228;
assign RESULT_u814=simplePinWrite_u232;
assign RESULT_u815=simplePinWrite_u229;
assign RESULT_u816=simplePinWrite_u231;
assign RESULT_u817=simplePinWrite;
assign RESULT_u818=simplePinWrite_u230;
assign DONE=reg_4fbb82fa_result_delayed_u0;
endmodule



module image1_iunzip_stateVar_In1PortEnable(bus_6b4f1791_, bus_7b3d8b32_, bus_1712d9e1_, bus_1301d8aa_, bus_71ee2f20_);
input		bus_6b4f1791_;
input		bus_7b3d8b32_;
input		bus_1712d9e1_;
input		bus_1301d8aa_;
output		bus_71ee2f20_;
reg		stateVar_In1PortEnable_u0=1'h0;
assign bus_71ee2f20_=stateVar_In1PortEnable_u0;
always @(posedge bus_6b4f1791_ or posedge bus_7b3d8b32_)
begin
if (bus_7b3d8b32_)
stateVar_In1PortEnable_u0<=1'h0;
else if (bus_1712d9e1_)
stateVar_In1PortEnable_u0<=bus_1301d8aa_;
end
endmodule



module image1_iunzip_firstNPixels(CLK, RESET, GO, port_0e7ec45d_, port_10601e70_, port_328b25f5_, port_33fbecb1_, port_30f2a2a5_, port_58472f4a_, RESULT, RESULT_u819, RESULT_u820, RESULT_u821, RESULT_u822, RESULT_u823, RESULT_u824, RESULT_u825, RESULT_u826, RESULT_u827, RESULT_u828, RESULT_u829, DONE);
input		CLK;
input		RESET;
input		GO;
input	[31:0]	port_0e7ec45d_;
input		port_10601e70_;
input		port_328b25f5_;
input	[15:0]	port_33fbecb1_;
input		port_30f2a2a5_;
input	[15:0]	port_58472f4a_;
output		RESULT;
output	[31:0]	RESULT_u819;
output		RESULT_u820;
output	[31:0]	RESULT_u821;
output	[15:0]	RESULT_u822;
output	[2:0]	RESULT_u823;
output		RESULT_u824;
output	[31:0]	RESULT_u825;
output	[2:0]	RESULT_u826;
output		RESULT_u827;
output	[31:0]	RESULT_u828;
output	[2:0]	RESULT_u829;
output		DONE;
wire		and_u1412_u0;
wire		and_u1413_u0;
wire	[31:0]	add;
wire		and_u1414_u0;
wire		or_u378_u0;
reg		reg_4854b0ab_u0=1'h0;
wire		or_u379_u0;
wire		and_u1415_u0;
reg		reg_4e678d3d_u0=1'h0;
reg	[15:0]	syncEnable_u99=16'h0;
reg		reg_72b58ef9_u0=1'h0;
reg		reg_72b58ef9_result_delayed_u0=1'h0;
reg		reg_4fa2b10d_u0=1'h0;
reg	[15:0]	syncEnable_u100_u0=16'h0;
wire	[15:0]	mux_u111;
wire		or_u380_u0;
wire	[31:0]	mux_u112_u0;
assign and_u1412_u0=GO&port_30f2a2a5_;
assign and_u1413_u0=GO&port_328b25f5_;
assign add=port_0e7ec45d_+32'h2;
assign and_u1414_u0=reg_4854b0ab_u0&port_10601e70_;
assign or_u378_u0=and_u1414_u0|RESET;
always @(posedge CLK or posedge reg_4fa2b10d_u0 or posedge or_u378_u0)
begin
if (or_u378_u0)
reg_4854b0ab_u0<=1'h0;
else if (reg_4fa2b10d_u0)
reg_4854b0ab_u0<=1'h1;
else reg_4854b0ab_u0<=reg_4854b0ab_u0;
end
assign or_u379_u0=and_u1415_u0|RESET;
assign and_u1415_u0=reg_4e678d3d_u0&port_10601e70_;
always @(posedge CLK or posedge reg_72b58ef9_u0 or posedge or_u379_u0)
begin
if (or_u379_u0)
reg_4e678d3d_u0<=1'h0;
else if (reg_72b58ef9_u0)
reg_4e678d3d_u0<=1'h1;
else reg_4e678d3d_u0<=reg_4e678d3d_u0;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u99<=port_33fbecb1_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_72b58ef9_u0<=1'h0;
else reg_72b58ef9_u0<=reg_4fa2b10d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_72b58ef9_result_delayed_u0<=1'h0;
else reg_72b58ef9_result_delayed_u0<=reg_72b58ef9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4fa2b10d_u0<=1'h0;
else reg_4fa2b10d_u0<=GO;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u100_u0<=port_58472f4a_;
end
assign mux_u111=(reg_4fa2b10d_u0)?syncEnable_u100_u0:syncEnable_u99;
assign or_u380_u0=reg_4fa2b10d_u0|reg_72b58ef9_u0;
assign mux_u112_u0=(reg_4fa2b10d_u0)?32'h0:32'h1;
assign RESULT=GO;
assign RESULT_u819=add;
assign RESULT_u820=or_u380_u0;
assign RESULT_u821={31'b0, mux_u112_u0[0]};
assign RESULT_u822=mux_u111;
assign RESULT_u823=3'h1;
assign RESULT_u824=GO;
assign RESULT_u825=32'h1;
assign RESULT_u826=3'h1;
assign RESULT_u827=GO;
assign RESULT_u828=32'h0;
assign RESULT_u829=3'h1;
assign DONE=reg_72b58ef9_result_delayed_u0;
endmodule



module image1_iunzip_simplememoryreferee_12559ca8_(bus_34d6401e_, bus_2c677a40_, bus_61602789_, bus_520a81dd_, bus_4f242077_, bus_56e7637f_, bus_2414a2f1_, bus_4906a1e5_, bus_0cb5957a_, bus_4c5426bf_, bus_4034cf94_, bus_12ed058a_, bus_50e7e991_, bus_4f572e1e_, bus_20b4c307_, bus_32b5a413_, bus_4b85717f_, bus_3181df50_, bus_2f2a289d_, bus_25006614_, bus_4d322080_, bus_77aca28c_, bus_6af53624_, bus_0a775a74_, bus_628ee2f9_, bus_0d379228_, bus_1e395c9f_, bus_3b62cf1f_, bus_4b0b58ac_, bus_6b5b6b3c_, bus_3c871d5b_, bus_225c3717_, bus_0cf04c6c_, bus_05e31049_, bus_32560469_, bus_1066ab06_, bus_52b719e4_, bus_08315480_);
input		bus_34d6401e_;
input		bus_2c677a40_;
input		bus_61602789_;
input	[15:0]	bus_520a81dd_;
input		bus_4f242077_;
input	[15:0]	bus_56e7637f_;
input	[31:0]	bus_2414a2f1_;
input	[2:0]	bus_4906a1e5_;
input		bus_0cb5957a_;
input		bus_4c5426bf_;
input	[15:0]	bus_4034cf94_;
input	[31:0]	bus_12ed058a_;
input	[2:0]	bus_50e7e991_;
input		bus_4f572e1e_;
input		bus_20b4c307_;
input	[15:0]	bus_32b5a413_;
input	[31:0]	bus_4b85717f_;
input	[2:0]	bus_3181df50_;
input		bus_2f2a289d_;
input	[31:0]	bus_25006614_;
input	[2:0]	bus_4d322080_;
input		bus_77aca28c_;
input	[31:0]	bus_6af53624_;
input	[2:0]	bus_0a775a74_;
output	[15:0]	bus_628ee2f9_;
output	[31:0]	bus_0d379228_;
output		bus_1e395c9f_;
output		bus_3b62cf1f_;
output	[2:0]	bus_4b0b58ac_;
output		bus_6b5b6b3c_;
output	[15:0]	bus_3c871d5b_;
output		bus_225c3717_;
output	[15:0]	bus_0cf04c6c_;
output		bus_05e31049_;
output	[15:0]	bus_32560469_;
output		bus_1066ab06_;
output	[15:0]	bus_52b719e4_;
output		bus_08315480_;
wire		or_35e97769_u0;
wire		or_2a51fa90_u0;
wire		not_1d76be37_u0;
wire		or_55542316_u0;
wire		and_21ff797d_u0;
wire		not_356cbbe8_u0;
wire		not_3e60f7a5_u0;
wire		or_46b4d4e4_u0;
wire		not_6a30a1a5_u0;
wire		or_2ee69eb0_u0;
wire	[15:0]	mux_703fee27_u0;
wire		or_12ad4cb5_u0;
reg		done_qual_u48_u0=1'h0;
wire	[31:0]	mux_34e90777_u0;
wire		and_45367429_u0;
reg		done_qual_u49_u0=1'h0;
wire		and_10c38621_u0;
wire		and_464ccae5_u0;
wire		not_6093bfb9_u0;
wire		or_12140f39_u0;
reg		done_qual_u50_u0=1'h0;
wire		or_7a84c33d_u0;
wire		and_771baaa0_u0;
reg		done_qual_u51_u0=1'h0;
wire		or_1968ad54_u0;
reg		done_qual_u52_u0=1'h0;
assign or_35e97769_u0=or_12140f39_u0|done_qual_u49_u0;
assign or_2a51fa90_u0=bus_4f242077_|done_qual_u52_u0;
assign not_1d76be37_u0=~bus_61602789_;
assign or_55542316_u0=bus_0cb5957a_|bus_4c5426bf_;
assign and_21ff797d_u0=or_35e97769_u0&bus_61602789_;
assign not_356cbbe8_u0=~bus_61602789_;
assign not_3e60f7a5_u0=~bus_61602789_;
assign or_46b4d4e4_u0=bus_77aca28c_|done_qual_u51_u0;
assign not_6a30a1a5_u0=~bus_61602789_;
assign or_2ee69eb0_u0=bus_4f242077_|bus_4c5426bf_|bus_20b4c307_;
assign mux_703fee27_u0=({16{bus_4f242077_}}&bus_56e7637f_)|({16{bus_4c5426bf_}}&bus_4034cf94_)|({16{bus_20b4c307_}}&bus_32b5a413_);
assign or_12ad4cb5_u0=bus_2f2a289d_|done_qual_u48_u0;
always @(posedge bus_34d6401e_)
begin
if (bus_2c677a40_)
done_qual_u48_u0<=1'h0;
else done_qual_u48_u0<=bus_2f2a289d_;
end
assign mux_34e90777_u0=({32{bus_4f242077_}}&{31'b0, bus_2414a2f1_[0]})|({32{or_55542316_u0}}&bus_12ed058a_)|({32{or_12140f39_u0}}&bus_4b85717f_)|({32{bus_2f2a289d_}}&bus_25006614_)|({32{bus_77aca28c_}}&bus_6af53624_);
assign and_45367429_u0=or_46b4d4e4_u0&bus_61602789_;
always @(posedge bus_34d6401e_)
begin
if (bus_2c677a40_)
done_qual_u49_u0<=1'h0;
else done_qual_u49_u0<=or_12140f39_u0;
end
assign and_10c38621_u0=or_12ad4cb5_u0&bus_61602789_;
assign bus_628ee2f9_=mux_703fee27_u0;
assign bus_0d379228_=mux_34e90777_u0;
assign bus_1e395c9f_=or_2ee69eb0_u0;
assign bus_3b62cf1f_=or_7a84c33d_u0;
assign bus_4b0b58ac_=3'h1;
assign bus_6b5b6b3c_=and_771baaa0_u0;
assign bus_3c871d5b_=bus_520a81dd_;
assign bus_225c3717_=and_464ccae5_u0;
assign bus_0cf04c6c_=bus_520a81dd_;
assign bus_05e31049_=and_21ff797d_u0;
assign bus_32560469_=bus_520a81dd_;
assign bus_1066ab06_=and_10c38621_u0;
assign bus_52b719e4_=bus_520a81dd_;
assign bus_08315480_=and_45367429_u0;
assign and_464ccae5_u0=or_1968ad54_u0&bus_61602789_;
assign not_6093bfb9_u0=~bus_61602789_;
assign or_12140f39_u0=bus_4f572e1e_|bus_20b4c307_;
always @(posedge bus_34d6401e_)
begin
if (bus_2c677a40_)
done_qual_u50_u0<=1'h0;
else done_qual_u50_u0<=or_55542316_u0;
end
assign or_7a84c33d_u0=bus_4f242077_|or_55542316_u0|or_12140f39_u0|bus_2f2a289d_|bus_77aca28c_;
assign and_771baaa0_u0=or_2a51fa90_u0&bus_61602789_;
always @(posedge bus_34d6401e_)
begin
if (bus_2c677a40_)
done_qual_u51_u0<=1'h0;
else done_qual_u51_u0<=bus_77aca28c_;
end
assign or_1968ad54_u0=or_55542316_u0|done_qual_u50_u0;
always @(posedge bus_34d6401e_)
begin
if (bus_2c677a40_)
done_qual_u52_u0<=1'h0;
else done_qual_u52_u0<=bus_4f242077_;
end
endmodule


