// __  ___ __ ___  _ __   ___  ___ 
// \ \/ / '__/ _ \| '_ \ / _ \/ __|
//  >  <| | | (_) | | | | (_) \__ \
// /_/\_\_|  \___/|_| |_|\___/|___/
// 
// Xronos synthesizer version
// Run date: Thu 2 Nov 2017 13:58:52 +0000
// 

module resized_HH2_xy(Out1_RDY, Out1_SEND, In1_ACK, Out1_COUNT, RESET, In1_SEND, In1_DATA, CLK, Out1_ACK, In1_COUNT, Out1_DATA);
input		Out1_RDY;
wire		consumeRow_done;
output		Out1_SEND;
wire		reset_go;
output		In1_ACK;
output	[15:0]	Out1_COUNT;
input		RESET;
input		In1_SEND;
input	[15:0]	In1_DATA;
wire		repeatRowExpanded_done;
input		CLK;
wire		consumeRow_go;
input		Out1_ACK;
wire		repeatRowExpanded_go;
wire		reset_done;
input	[15:0]	In1_COUNT;
output	[15:0]	Out1_DATA;
wire		bus_5c918e28_;
wire		bus_24921465_;
wire	[15:0]	scheduler_u217;
wire	[15:0]	scheduler_u216;
wire		resized_HH2_xy_scheduler_instance_DONE;
wire		scheduler_u207;
wire		scheduler_u214;
wire	[31:0]	scheduler_u200;
wire	[31:0]	scheduler_u204;
wire	[31:0]	scheduler_u206;
wire	[31:0]	scheduler_u210;
wire		scheduler_u205;
wire		scheduler;
wire	[2:0]	scheduler_u211;
wire		scheduler_u203;
wire		scheduler_u201;
wire		scheduler_u212;
wire		scheduler_u215;
wire		scheduler_u202;
wire		scheduler_u208;
wire		scheduler_u209;
wire		scheduler_u213;
wire	[31:0]	bus_159d7a35_;
wire	[15:0]	bus_084c0cb4_;
wire		bus_749f2f87_;
wire		bus_2635a5e4_;
wire		bus_68a9d0f3_;
wire	[15:0]	bus_046d1002_;
wire		bus_6a6e976a_;
wire	[15:0]	bus_3fd024dd_;
wire	[31:0]	bus_0b94f26f_;
wire		bus_6390af6d_;
wire	[15:0]	bus_5931117b_;
wire	[31:0]	bus_2ae1483e_;
wire	[15:0]	bus_7a3d3bb9_;
wire	[31:0]	bus_46701177_;
wire		bus_37b58ffd_;
wire		bus_6ae64912_;
wire	[2:0]	bus_43e739c0_;
wire		bus_70595e48_;
wire		bus_1caadeaa_;
wire	[15:0]	bus_7faadc73_;
wire		bus_480a5dc4_;
wire	[31:0]	consumeRow_u16;
wire	[2:0]	consumeRow_u14;
wire	[2:0]	consumeRow_u18;
wire	[31:0]	consumeRow_u12;
wire		consumeRow_u15;
wire	[15:0]	consumeRow_u17;
wire		consumeRow_u11;
wire		resized_HH2_xy_consumeRow_instance_DONE;
wire		consumeRow;
wire	[15:0]	consumeRow_u10;
wire		consumeRow_u19;
wire	[15:0]	consumeRow_u13;
wire	[31:0]	repeatRowExpanded_u13;
wire	[15:0]	repeatRowExpanded_u14;
wire	[15:0]	repeatRowExpanded_u8;
wire		repeatRowExpanded_u9;
wire		resized_HH2_xy_repeatRowExpanded_instance_DONE;
wire		repeatRowExpanded_u12;
wire	[2:0]	repeatRowExpanded_u11;
wire		repeatRowExpanded;
wire	[31:0]	repeatRowExpanded_u10;
wire	[2:0]	repeatRowExpanded_u15;
wire		bus_59c83a2c_;
wire		bus_0b61c797_;
wire	[2:0]	bus_13e0228b_;
wire		bus_1b9989aa_;
wire		bus_15d988f3_;
wire	[15:0]	bus_08f43ee3_;
wire	[15:0]	bus_27c6803d_;
wire		bus_7fa5bd8d_;
wire	[31:0]	bus_5fed9ad9_;
wire		bus_2570462b_;
wire		reset;
wire		reset_u4;
wire	[15:0]	reset_u3;
wire	[15:0]	reset_u5;
wire		resized_HH2_xy_reset_instance_DONE;
assign consumeRow_done=bus_24921465_;
assign Out1_SEND=scheduler_u213;
assign reset_go=scheduler_u215;
assign In1_ACK=consumeRow_u19;
assign Out1_COUNT=scheduler_u216;
assign repeatRowExpanded_done=bus_6390af6d_;
assign consumeRow_go=scheduler_u212;
assign repeatRowExpanded_go=scheduler_u214;
assign reset_done=bus_59c83a2c_;
assign Out1_DATA=scheduler_u217;
resized_HH2_xy_Kicker_39 resized_HH2_xy_Kicker_39_1(.CLK(CLK), .RESET(bus_0b61c797_), 
  .bus_5c918e28_(bus_5c918e28_));
assign bus_24921465_=resized_HH2_xy_consumeRow_instance_DONE&{1{resized_HH2_xy_consumeRow_instance_DONE}};
resized_HH2_xy_scheduler resized_HH2_xy_scheduler_instance(.CLK(CLK), .RESET(bus_0b61c797_), 
  .GO(bus_5c918e28_), .port_4e51436e_(32'h0), .port_768be70f_(bus_6a6e976a_), .port_30496c3f_(bus_159d7a35_), 
  .port_1bf015b7_(bus_0b94f26f_), .port_607140ed_(bus_2635a5e4_), .port_038b3c60_(bus_5931117b_), 
  .port_7451eb09_(bus_3fd024dd_), .port_4a47b2ff_(bus_6ae64912_), .port_7dc406cd_(bus_7faadc73_), 
  .port_6a29d19a_(Out1_RDY), .port_19608f97_(consumeRow_done), .port_1372f033_(reset_done), 
  .port_32809d55_(repeatRowExpanded_done), .port_1bbb1093_(In1_SEND), .DONE(resized_HH2_xy_scheduler_instance_DONE), 
  .RESULT(scheduler), .RESULT_u1334(scheduler_u200), .RESULT_u1335(scheduler_u201), 
  .RESULT_u1336(scheduler_u202), .RESULT_u1337(scheduler_u203), .RESULT_u1338(scheduler_u204), 
  .RESULT_u1339(scheduler_u205), .RESULT_u1340(scheduler_u206), .RESULT_u1341(scheduler_u207), 
  .RESULT_u1342(scheduler_u208), .RESULT_u1343(scheduler_u209), .RESULT_u1344(scheduler_u210), 
  .RESULT_u1345(scheduler_u211), .RESULT_u1346(scheduler_u212), .RESULT_u1347(scheduler_u213), 
  .RESULT_u1348(scheduler_u214), .RESULT_u1349(scheduler_u215), .RESULT_u1350(scheduler_u216), 
  .RESULT_u1351(scheduler_u217));
resized_HH2_xy_stateVar_Out1TokenIndex resized_HH2_xy_stateVar_Out1TokenIndex_1(.bus_7ed6fa76_(CLK), 
  .bus_763548e3_(bus_0b61c797_), .bus_51456afc_(scheduler_u203), .bus_44270e5a_(scheduler_u204), 
  .bus_159d7a35_(bus_159d7a35_));
resized_HH2_xy_structuralmemory_2116ed52_ resized_HH2_xy_structuralmemory_2116ed52__1(.CLK_u11(CLK), 
  .bus_3407a066_(bus_0b61c797_), .bus_02a6eccb_(bus_5fed9ad9_), .bus_404a7c0c_(3'h1), 
  .bus_7ff7fda2_(bus_2570462b_), .bus_05f7b94c_(bus_1b9989aa_), .bus_5ba84a22_(bus_27c6803d_), 
  .bus_084c0cb4_(bus_084c0cb4_), .bus_749f2f87_(bus_749f2f87_));
resized_HH2_xy_stateVar_Out1PortEnable resized_HH2_xy_stateVar_Out1PortEnable_1(.bus_6395a33f_(CLK), 
  .bus_160e9142_(bus_0b61c797_), .bus_4d5774e5_(scheduler_u207), .bus_6173af9a_(scheduler_u208), 
  .bus_2635a5e4_(bus_2635a5e4_));
resized_HH2_xy_structuralmemory_121950d1_ resized_HH2_xy_structuralmemory_121950d1__1(.CLK_u12(CLK), 
  .bus_1b9eeab7_(bus_0b61c797_), .bus_4a6c0845_(bus_46701177_), .bus_0355a864_(3'h1), 
  .bus_00c34d18_(bus_480a5dc4_), .bus_200222a1_(bus_1caadeaa_), .bus_4aa3f2c6_(bus_7a3d3bb9_), 
  .bus_046d1002_(bus_046d1002_), .bus_68a9d0f3_(bus_68a9d0f3_));
resized_HH2_xy_stateVar_fsmState_resized_HH2_xy resized_HH2_xy_stateVar_fsmState_resized_HH2_xy_1(.bus_027c1c08_(CLK), 
  .bus_1040e6d7_(bus_0b61c797_), .bus_1c5da006_(scheduler_u201), .bus_69c25494_(scheduler_u202), 
  .bus_6a6e976a_(bus_6a6e976a_));
resized_HH2_xy_stateVar_rowRepeated resized_HH2_xy_stateVar_rowRepeated_1(.bus_49b93211_(CLK), 
  .bus_0c3dac10_(bus_0b61c797_), .bus_58b6be80_(repeatRowExpanded), .bus_39234c02_(repeatRowExpanded_u8), 
  .bus_4e9c8a8a_(reset), .bus_4cf3f116_(16'h1), .bus_3fd024dd_(bus_3fd024dd_));
resized_HH2_xy_stateVar_Out1MaxTokenIndex resized_HH2_xy_stateVar_Out1MaxTokenIndex_1(.bus_2fb5cc44_(CLK), 
  .bus_2eaa1fa7_(bus_0b61c797_), .bus_0662c425_(scheduler_u205), .bus_799d8f37_(scheduler_u206), 
  .bus_0b94f26f_(bus_0b94f26f_));
assign bus_6390af6d_=resized_HH2_xy_repeatRowExpanded_instance_DONE&{1{resized_HH2_xy_repeatRowExpanded_instance_DONE}};
resized_HH2_xy_stateVar_x resized_HH2_xy_stateVar_x_1(.bus_2e51ce68_(CLK), .bus_365ac0ca_(bus_0b61c797_), 
  .bus_5f0f6c4a_(consumeRow), .bus_1f3118e6_(consumeRow_u10), .bus_2341ca1a_(reset_u4), 
  .bus_25e6f202_(16'h0), .bus_5931117b_(bus_5931117b_));
resized_HH2_xy_stateVar_fsmOldState_resized_HH2_xy resized_HH2_xy_stateVar_fsmOldState_resized_HH2_xy_1(.bus_5900bf5a_(CLK), 
  .bus_353bfc63_(bus_0b61c797_), .bus_58660ccc_(scheduler), .bus_6ef2aeea_(32'h0), 
  .bus_2ae1483e_(bus_2ae1483e_));
resized_HH2_xy_simplememoryreferee_390f3e2f_ resized_HH2_xy_simplememoryreferee_390f3e2f__1(.bus_23993a97_(CLK), 
  .bus_7cef1f98_(bus_0b61c797_), .bus_7ebc765f_(bus_68a9d0f3_), .bus_2d8c8d97_(bus_046d1002_), 
  .bus_71cc810b_(consumeRow_u15), .bus_7a8a14d8_(consumeRow_u17), .bus_706609c9_(consumeRow_u16), 
  .bus_2df6d93b_(3'h1), .bus_2ded108e_(repeatRowExpanded_u12), .bus_2e3a2c30_(repeatRowExpanded_u14), 
  .bus_14e3e00d_(repeatRowExpanded_u13), .bus_194afe2d_(3'h1), .bus_647b7d66_(scheduler_u209), 
  .bus_4b65d917_(scheduler_u210), .bus_4edd6dce_(3'h1), .bus_7a3d3bb9_(bus_7a3d3bb9_), 
  .bus_46701177_(bus_46701177_), .bus_1caadeaa_(bus_1caadeaa_), .bus_480a5dc4_(bus_480a5dc4_), 
  .bus_43e739c0_(bus_43e739c0_), .bus_70595e48_(bus_70595e48_), .bus_37b58ffd_(bus_37b58ffd_), 
  .bus_7faadc73_(bus_7faadc73_), .bus_6ae64912_(bus_6ae64912_));
resized_HH2_xy_consumeRow resized_HH2_xy_consumeRow_instance(.CLK(CLK), .RESET(bus_0b61c797_), 
  .GO(consumeRow_go), .port_0bc8ac8b_(bus_5931117b_), .port_3de2b1d0_(bus_15d988f3_), 
  .port_01480d6c_(bus_70595e48_), .port_43c4e7d2_(In1_DATA), .DONE(resized_HH2_xy_consumeRow_instance_DONE), 
  .RESULT(consumeRow), .RESULT_u1352(consumeRow_u10), .RESULT_u1353(consumeRow_u11), 
  .RESULT_u1354(consumeRow_u12), .RESULT_u1355(consumeRow_u13), .RESULT_u1356(consumeRow_u14), 
  .RESULT_u1357(consumeRow_u15), .RESULT_u1358(consumeRow_u16), .RESULT_u1359(consumeRow_u17), 
  .RESULT_u1360(consumeRow_u18), .RESULT_u1361(consumeRow_u19));
resized_HH2_xy_repeatRowExpanded resized_HH2_xy_repeatRowExpanded_instance(.CLK(CLK), 
  .RESET(bus_0b61c797_), .GO(repeatRowExpanded_go), .port_3ddff29c_(bus_3fd024dd_), 
  .port_42abce2f_(bus_7fa5bd8d_), .port_6af401d3_(bus_08f43ee3_), .port_516974d5_(bus_37b58ffd_), 
  .DONE(resized_HH2_xy_repeatRowExpanded_instance_DONE), .RESULT(repeatRowExpanded), 
  .RESULT_u1362(repeatRowExpanded_u8), .RESULT_u1363(repeatRowExpanded_u9), .RESULT_u1364(repeatRowExpanded_u10), 
  .RESULT_u1365(repeatRowExpanded_u11), .RESULT_u1366(repeatRowExpanded_u12), 
  .RESULT_u1367(repeatRowExpanded_u13), .RESULT_u1368(repeatRowExpanded_u14), 
  .RESULT_u1369(repeatRowExpanded_u15));
assign bus_59c83a2c_=resized_HH2_xy_reset_instance_DONE&{1{resized_HH2_xy_reset_instance_DONE}};
resized_HH2_xy_globalreset_physical_08a74754_ resized_HH2_xy_globalreset_physical_08a74754__1(.bus_139efad7_(CLK), 
  .bus_67634e72_(RESET), .bus_0b61c797_(bus_0b61c797_));
resized_HH2_xy_simplememoryreferee_519aba6e_ resized_HH2_xy_simplememoryreferee_519aba6e__1(.bus_31e46996_(CLK), 
  .bus_78041c94_(bus_0b61c797_), .bus_69efc929_(bus_749f2f87_), .bus_09bbc993_(bus_084c0cb4_), 
  .bus_3ec76267_(consumeRow_u11), .bus_4f50e209_(consumeRow_u13), .bus_3cbefa4e_(consumeRow_u12), 
  .bus_57eee443_(3'h1), .bus_5133aa26_(repeatRowExpanded_u9), .bus_649a3ec9_(repeatRowExpanded_u10), 
  .bus_7184d705_(3'h1), .bus_27c6803d_(bus_27c6803d_), .bus_5fed9ad9_(bus_5fed9ad9_), 
  .bus_1b9989aa_(bus_1b9989aa_), .bus_2570462b_(bus_2570462b_), .bus_13e0228b_(bus_13e0228b_), 
  .bus_15d988f3_(bus_15d988f3_), .bus_08f43ee3_(bus_08f43ee3_), .bus_7fa5bd8d_(bus_7fa5bd8d_));
resized_HH2_xy_reset resized_HH2_xy_reset_instance(.CLK(CLK), .RESET(bus_0b61c797_), 
  .GO(reset_go), .DONE(resized_HH2_xy_reset_instance_DONE), .RESULT(reset), .RESULT_u1370(reset_u3), 
  .RESULT_u1371(reset_u4), .RESULT_u1372(reset_u5));
endmodule



module resized_HH2_xy_Kicker_39(CLK, RESET, bus_5c918e28_);
input		CLK;
input		RESET;
output		bus_5c918e28_;
wire		bus_6a1c8991_;
reg		kicker_2=1'h0;
wire		bus_7e97e12a_;
reg		kicker_res=1'h0;
wire		bus_1fbd5a84_;
reg		kicker_1=1'h0;
wire		bus_7c192699_;
assign bus_6a1c8991_=bus_7e97e12a_&kicker_1;
always @(posedge CLK)
begin
kicker_2<=bus_6a1c8991_;
end
assign bus_7e97e12a_=~RESET;
always @(posedge CLK)
begin
kicker_res<=bus_7c192699_;
end
assign bus_5c918e28_=kicker_res;
assign bus_1fbd5a84_=~kicker_2;
always @(posedge CLK)
begin
kicker_1<=bus_7e97e12a_;
end
assign bus_7c192699_=kicker_1&bus_7e97e12a_&bus_1fbd5a84_;
endmodule



module resized_HH2_xy_scheduler(CLK, RESET, GO, port_4e51436e_, port_768be70f_, port_30496c3f_, port_1bf015b7_, port_607140ed_, port_038b3c60_, port_7451eb09_, port_4a47b2ff_, port_7dc406cd_, port_6a29d19a_, port_19608f97_, port_1372f033_, port_32809d55_, port_1bbb1093_, RESULT, RESULT_u1334, RESULT_u1335, RESULT_u1336, RESULT_u1337, RESULT_u1338, RESULT_u1339, RESULT_u1340, RESULT_u1341, RESULT_u1342, RESULT_u1343, RESULT_u1344, RESULT_u1345, RESULT_u1346, RESULT_u1347, RESULT_u1348, RESULT_u1349, RESULT_u1350, RESULT_u1351, DONE);
input		CLK;
input		RESET;
input		GO;
input	[31:0]	port_4e51436e_;
input		port_768be70f_;
input	[31:0]	port_30496c3f_;
input	[31:0]	port_1bf015b7_;
input		port_607140ed_;
input	[15:0]	port_038b3c60_;
input	[15:0]	port_7451eb09_;
input		port_4a47b2ff_;
input	[15:0]	port_7dc406cd_;
input		port_6a29d19a_;
input		port_19608f97_;
input		port_1372f033_;
input		port_32809d55_;
input		port_1bbb1093_;
output		RESULT;
output	[31:0]	RESULT_u1334;
output		RESULT_u1335;
output		RESULT_u1336;
output		RESULT_u1337;
output	[31:0]	RESULT_u1338;
output		RESULT_u1339;
output	[31:0]	RESULT_u1340;
output		RESULT_u1341;
output		RESULT_u1342;
output		RESULT_u1343;
output	[31:0]	RESULT_u1344;
output	[2:0]	RESULT_u1345;
output		RESULT_u1346;
output		RESULT_u1347;
output		RESULT_u1348;
output		RESULT_u1349;
output	[15:0]	RESULT_u1350;
output	[15:0]	RESULT_u1351;
output		DONE;
wire		lessThan;
wire	[15:0]	lessThan_a_unsigned;
wire	[15:0]	lessThan_b_unsigned;
wire	[15:0]	equals_a_unsigned;
wire		equals;
wire	[15:0]	equals_b_unsigned;
wire	[15:0]	lessThan_u50_b_unsigned;
wire	[15:0]	lessThan_u50_a_unsigned;
wire		lessThan_u50;
wire		andOp;
wire		equals_u116;
wire	[15:0]	equals_u116_a_unsigned;
wire	[15:0]	equals_u116_b_unsigned;
wire signed	[31:0]	equals_u117_b_signed;
wire		equals_u117;
wire signed	[31:0]	equals_u117_a_signed;
wire		and_u2210_u0;
wire		not_u405_u0;
wire		and_u2211_u0;
wire		andOp_u133;
wire		not_u406_u0;
wire		and_u2212_u0;
wire		and_u2213_u0;
wire		simplePinWrite;
wire		not_u407_u0;
wire		and_u2214_u0;
wire		and_u2215_u0;
wire		simplePinWrite_u366;
wire		and_u2216_u0;
wire		not_u408_u0;
wire		and_u2217_u0;
wire		simplePinWrite_u367;
wire		and_u2218_u0;
reg		reg_62bcd2be_u0=1'h0;
reg		reg_64049807_u0=1'h0;
reg		reg_5c7b4c7d_u0=1'h0;
reg		reg_1cd8b4df_u0=1'h0;
reg		reg_640dac03_u0=1'h0;
reg		reg_7e3e122c_u0=1'h0;
reg		reg_0b38372d_u0=1'h0;
reg		reg_710efd1b_u0=1'h0;
reg		reg_2a321227_u0=1'h0;
reg		reg_36ce22d8_u0=1'h0;
reg		reg_6bf613ee_u0=1'h0;
reg		reg_18ad0cb7_u0=1'h0;
reg		reg_30e4f8f8_u0=1'h0;
reg		reg_24a21cbf_u0=1'h0;
reg		reg_64daf8c4_u0=1'h0;
reg		reg_54ef10cf_u0=1'h0;
reg		reg_77668746_u0=1'h0;
reg		reg_77668746_result_delayed_u0=1'h0;
reg		reg_66565274_u0=1'h0;
reg		reg_6d759d56_u0=1'h0;
reg		reg_7bd0a7f4_u0=1'h0;
reg		reg_201eb03b_u0=1'h0;
reg		reg_7d231906_u0=1'h0;
reg		reg_42b58a90_u0=1'h0;
reg		reg_382aec0c_u0=1'h0;
reg		reg_1457ec7b_u0=1'h0;
reg		reg_02369e1a_u0=1'h0;
reg		reg_6848807a_u0=1'h0;
reg		reg_1a837eb0_u0=1'h0;
reg		reg_45a11597_u0=1'h0;
reg		reg_774ab77d_u0=1'h0;
reg		reg_62921ea8_u0=1'h0;
reg		reg_0034740f_u0=1'h0;
reg		reg_1a0fb632_u0=1'h0;
reg		reg_061a1224_u0=1'h0;
reg		reg_58a2a0e3_u0=1'h0;
reg		reg_027e723d_u0=1'h0;
reg		reg_39d6e99f_u0=1'h0;
reg		reg_576a3720_u0=1'h0;
reg		reg_30e4f8f8_result_delayed_u0=1'h0;
reg		reg_00af20e1_u0=1'h0;
reg		reg_532c937d_u0=1'h0;
reg		reg_228ef2dc_u0=1'h0;
reg		reg_02369e1a_result_delayed_u0=1'h0;
reg		reg_0d9b29cf_u0=1'h0;
reg		reg_1098e4cf_u0=1'h0;
reg		reg_47aed7f7_u0=1'h0;
reg		reg_0ced50b0_u0=1'h0;
reg		reg_6d17e172_u0=1'h0;
reg		reg_75fb999e_u0=1'h0;
reg		reg_5046f020_u0=1'h0;
reg		reg_579a33fd_u0=1'h0;
reg		reg_53090f63_u0=1'h0;
reg		reg_38a628ca_u0=1'h0;
reg		reg_6a79fa17_u0=1'h0;
reg		reg_02369e1a_result_delayed_result_delayed_u0=1'h0;
reg		reg_7d46a529_u0=1'h0;
reg		reg_06efce9a_u0=1'h0;
reg		reg_1a0fb632_result_delayed_u0=1'h0;
reg		reg_24a21cbf_result_delayed_u0=1'h0;
reg		reg_4cd00ca8_u0=1'h0;
reg		reg_39c815b1_u0=1'h0;
reg		reg_229d1ee4_u0=1'h0;
reg		reg_4cc74cbd_u0=1'h0;
reg		reg_6d923de9_u0=1'h0;
reg		reg_0b8053fe_u0=1'h0;
reg		reg_06dc9aa2_u0=1'h0;
reg		reg_796241e6_u0=1'h0;
reg		reg_0425c0a1_u0=1'h0;
reg		reg_4a77e6f2_u0=1'h0;
reg		reg_387904fe_u0=1'h0;
reg		reg_3c2e9ca2_u0=1'h0;
reg		reg_66c4e649_u0=1'h0;
reg		reg_010c659c_u0=1'h0;
reg		reg_774ab77d_result_delayed_u0=1'h0;
reg		reg_4cc74cbd_result_delayed_u0=1'h0;
reg		reg_1f1eb78a_u0=1'h0;
reg		reg_0346d3d3_u0=1'h0;
reg		reg_6a895611_u0=1'h0;
wire		and_u2219_u0;
reg		reg_242facb3_u0=1'h0;
reg		reg_747c90de_u0=1'h0;
reg		reg_38a0bc03_u0=1'h0;
reg		reg_31615dc2_u0=1'h0;
reg		reg_10810426_u0=1'h0;
reg		reg_7a05baae_u0=1'h0;
reg		reg_68ca4866_u0=1'h0;
reg		reg_6ec6926a_u0=1'h0;
reg		reg_343e0093_u0=1'h0;
reg		reg_0b8053fe_result_delayed_u0=1'h0;
reg		reg_0ee3ba53_u0=1'h0;
reg		reg_2894b025_u0=1'h0;
reg		reg_03b6ff07_u0=1'h0;
reg		reg_49242595_u0=1'h0;
reg		reg_1680ee34_u0=1'h0;
reg		reg_1dd4f561_u0=1'h0;
reg		reg_13b25f04_u0=1'h0;
reg		reg_06efce9a_result_delayed_u0=1'h0;
reg		reg_48ad5013_u0=1'h0;
reg		reg_1c7bd8c5_u0=1'h0;
reg		reg_31a64119_u0=1'h0;
reg		reg_0fa7db18_u0=1'h0;
reg		reg_2c1074d0_u0=1'h0;
reg		reg_09a32d61_u0=1'h0;
reg		reg_77d7ef15_u0=1'h0;
reg		reg_677157b7_u0=1'h0;
reg		reg_68e2082a_u0=1'h0;
reg		reg_29ad1d65_u0=1'h0;
reg		reg_6f2cfbe7_u0=1'h0;
reg		reg_34d4a805_u0=1'h0;
reg		reg_68801c52_u0=1'h0;
reg		reg_6092b844_u0=1'h0;
reg		reg_5ee7823f_u0=1'h0;
reg		reg_6d759d56_result_delayed_u0=1'h0;
reg		reg_35da3503_u0=1'h0;
reg		reg_4c9f1046_u0=1'h0;
reg		reg_142b80f2_u0=1'h0;
reg		reg_29984143_u0=1'h0;
reg		reg_1dff8122_u0=1'h0;
reg		reg_229d1ee4_result_delayed_u0=1'h0;
reg		reg_1dce6126_u0=1'h0;
reg		reg_6848807a_result_delayed_u0=1'h0;
reg		reg_42b58a90_result_delayed_u0=1'h0;
reg		reg_4a3f86cf_u0=1'h0;
reg		reg_5a7e368e_u0=1'h0;
reg		reg_62921ea8_result_delayed_u0=1'h0;
reg		reg_5bc0cf31_u0=1'h0;
reg		reg_6a895611_result_delayed_u0=1'h0;
reg		reg_62b86a49_u0=1'h0;
reg		reg_4589457b_u0=1'h0;
reg		reg_710f71fd_u0=1'h0;
reg		reg_6092b844_result_delayed_u0=1'h0;
reg		reg_6f2cfbe7_result_delayed_u0=1'h0;
reg		reg_1ea77ba6_u0=1'h0;
reg		reg_62921ea8_result_delayed_result_delayed_u0=1'h0;
reg		reg_24232921_u0=1'h0;
reg		reg_06dc9aa2_result_delayed_u0=1'h0;
reg		reg_33b2aabd_u0=1'h0;
reg		reg_5e4d335d_u0=1'h0;
reg		reg_38645974_u0=1'h0;
reg		reg_7010ad01_u0=1'h0;
reg		reg_0320d63a_u0=1'h0;
reg		reg_5e188306_u0=1'h0;
reg		reg_0fa7db18_result_delayed_u0=1'h0;
reg		reg_439b9ebb_u0=1'h0;
reg		reg_7d510c70_u0=1'h0;
reg		reg_367fcb5d_u0=1'h0;
reg		reg_4ec55fe6_u0=1'h0;
reg		reg_0ced50b0_result_delayed_u0=1'h0;
reg		reg_4e1c133b_u0=1'h0;
reg		reg_061a1224_result_delayed_u0=1'h0;
reg		reg_6092b844_result_delayed_result_delayed_u0=1'h0;
reg		reg_441fe928_u0=1'h0;
reg		reg_13cde2f7_u0=1'h0;
reg		reg_2d8f78b3_u0=1'h0;
reg		reg_4bbdc680_u0=1'h0;
reg		reg_258244c0_u0=1'h0;
reg		reg_06dc9aa2_result_delayed_result_delayed_u0=1'h0;
reg		reg_38a0bc03_result_delayed_u0=1'h0;
reg		reg_1418995e_u0=1'h0;
reg		reg_1036257e_u0=1'h0;
reg		reg_5e4d335d_result_delayed_u0=1'h0;
reg		reg_4a5adf10_u0=1'h0;
reg		reg_0f726638_u0=1'h0;
reg		reg_4ffb5ab4_u0=1'h0;
reg		reg_6848807a_result_delayed_result_delayed_u0=1'h0;
reg		reg_0f2ec27d_u0=1'h0;
reg		reg_35d48481_u0=1'h0;
reg		reg_6dec38b5_u0=1'h0;
reg		reg_5bc0cf31_result_delayed_u0=1'h0;
reg		reg_64049807_result_delayed_u0=1'h0;
reg		reg_04da25b8_u0=1'h0;
reg		reg_6320b243_u0=1'h0;
reg		reg_0a6a1b0e_u0=1'h0;
reg		reg_747c90de_result_delayed_u0=1'h0;
reg		reg_64e0b984_u0=1'h0;
reg		reg_42b58a90_result_delayed_result_delayed_u0=1'h0;
reg		reg_05b030d6_u0=1'h0;
reg		reg_4ca109c7_u0=1'h0;
reg		reg_3a15fb72_u0=1'h0;
reg		reg_55edd085_u0=1'h0;
reg		reg_0034740f_result_delayed_u0=1'h0;
reg		reg_6f9e56f4_u0=1'h0;
reg		reg_76ad5fc6_u0=1'h0;
reg		reg_6320b243_result_delayed_u0=1'h0;
reg		reg_1dd4f561_result_delayed_u0=1'h0;
reg		reg_0b38372d_result_delayed_u0=1'h0;
reg		reg_405c3132_u0=1'h0;
reg		reg_2ea3b7cc_u0=1'h0;
reg		reg_0076a506_u0=1'h0;
reg		reg_4a5adf10_result_delayed_u0=1'h0;
reg		reg_0b769204_u0=1'h0;
reg		reg_64789d0a_u0=1'h0;
reg		reg_56b4ebc1_u0=1'h0;
reg		reg_6c7e010b_u0=1'h0;
reg		reg_4ca109c7_result_delayed_u0=1'h0;
reg		reg_0cc8a5bf_u0=1'h0;
reg		reg_35da3503_result_delayed_u0=1'h0;
reg		reg_21c538b9_u0=1'h0;
reg		reg_6f9e56f4_result_delayed_u0=1'h0;
reg		reg_7ffc667d_u0=1'h0;
reg		reg_26133792_u0=1'h0;
reg		reg_4e289baa_u0=1'h0;
reg		reg_579a33fd_result_delayed_u0=1'h0;
reg		reg_710f71fd_result_delayed_u0=1'h0;
reg		reg_4cd00ca8_result_delayed_u0=1'h0;
reg		reg_382aec0c_result_delayed_u0=1'h0;
wire		or_u689_u0;
reg		reg_38a0bc03_result_delayed_result_delayed_u0=1'h0;
reg		reg_4e1c133b_result_delayed_u0=1'h0;
reg		reg_5674bffb_u0=1'h0;
reg		reg_4769eae6_u0=1'h0;
reg		reg_7a05baae_result_delayed_u0=1'h0;
reg		reg_3f8e0a19_u0=1'h0;
reg		reg_5c7b4c7d_result_delayed_u0=1'h0;
reg		reg_45a11597_result_delayed_u0=1'h0;
reg		reg_6c7e010b_result_delayed_u0=1'h0;
reg		reg_242facb3_result_delayed_u0=1'h0;
reg		reg_35c4a85b_u0=1'h0;
reg		reg_2efcd75c_u0=1'h0;
reg		reg_29984143_result_delayed_u0=1'h0;
reg		reg_6028598b_u0=1'h0;
reg		reg_0f5456f1_u0=1'h0;
reg		reg_28e37146_u0=1'h0;
reg		reg_42b58a90_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_77d7ef15_result_delayed_u0=1'h0;
reg		reg_4cd00ca8_result_delayed_result_delayed_u0=1'h0;
reg		reg_0986382d_u0=1'h0;
reg		reg_3ecadb64_u0=1'h0;
reg		reg_1a79d7d6_u0=1'h0;
reg		reg_22f13343_u0=1'h0;
reg		reg_32c8d37c_u0=1'h0;
reg		reg_4f367a8e_u0=1'h0;
reg		reg_76f5e34d_u0=1'h0;
reg		reg_0346d3d3_result_delayed_u0=1'h0;
reg		reg_7d212c9a_u0=1'h0;
reg		reg_64049807_result_delayed_result_delayed_u0=1'h0;
reg		reg_5101c4c6_u0=1'h0;
reg		reg_4589457b_result_delayed_u0=1'h0;
reg		reg_02369e1a_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_7a05baae_result_delayed_result_delayed_u0=1'h0;
reg		reg_42536b9e_u0=1'h0;
reg		reg_7010ad01_result_delayed_u0=1'h0;
reg		reg_40fef52d_u0=1'h0;
reg		reg_070292d1_u0=1'h0;
reg		reg_42b58a90_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_1c1149c7_u0=1'h0;
reg		reg_6028598b_result_delayed_u0=1'h0;
reg		reg_64049807_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_150760de_u0=1'h0;
reg		reg_104b8d92_u0=1'h0;
reg		reg_0ee3ba53_result_delayed_u0=1'h0;
reg		reg_7ffc667d_result_delayed_u0=1'h0;
reg		reg_38a628ca_result_delayed_u0=1'h0;
reg		reg_6df7e814_u0=1'h0;
reg		reg_5101c4c6_result_delayed_u0=1'h0;
reg		reg_1fa5ca42_u0=1'h0;
reg		reg_183f91d8_u0=1'h0;
reg		reg_2537f8df_u0=1'h0;
reg		reg_337b1691_u0=1'h0;
reg		reg_426d8380_u0=1'h0;
reg		reg_650388ee_u0=1'h0;
reg		reg_2894b025_result_delayed_u0=1'h0;
reg		reg_48ad5013_result_delayed_u0=1'h0;
reg		reg_68801c52_result_delayed_u0=1'h0;
reg		reg_09069cf0_u0=1'h0;
reg		reg_445ccdaa_u0=1'h0;
reg		reg_14de3123_u0=1'h0;
reg		reg_62bcd2be_result_delayed_u0=1'h0;
reg		reg_7338c2c5_u0=1'h0;
reg		reg_15c73839_u0=1'h0;
reg		reg_51172316_u0=1'h0;
reg		reg_1fbac5be_u0=1'h0;
reg		reg_4ffb5ab4_result_delayed_u0=1'h0;
reg		reg_5a7e368e_result_delayed_u0=1'h0;
reg		reg_38a628ca_result_delayed_result_delayed_u0=1'h0;
reg		reg_6f9e56f4_result_delayed_result_delayed_u0=1'h0;
reg		reg_75ddf3cd_u0=1'h0;
reg		reg_222ee43c_u0=1'h0;
reg		reg_24232921_result_delayed_u0=1'h0;
reg		reg_2a60e877_u0=1'h0;
reg		reg_1c7bd8c5_result_delayed_u0=1'h0;
reg		reg_05b030d6_result_delayed_u0=1'h0;
reg		reg_6df7e814_result_delayed_u0=1'h0;
reg		reg_0530331a_u0=1'h0;
reg		reg_5df79fda_u0=1'h0;
reg		reg_2add40ec_u0=1'h0;
reg		reg_195de36c_u0=1'h0;
reg		reg_4f367a8e_result_delayed_u0=1'h0;
reg		reg_70b8aa8a_u0=1'h0;
reg		reg_52bc0089_u0=1'h0;
reg		reg_0fa7db18_result_delayed_result_delayed_u0=1'h0;
reg		reg_62bcd2be_result_delayed_result_delayed_u0=1'h0;
reg		reg_01a00b9a_u0=1'h0;
reg		reg_08eb52d0_u0=1'h0;
reg		reg_68801c52_result_delayed_result_delayed_u0=1'h0;
reg		reg_66565274_result_delayed_u0=1'h0;
reg		reg_3c2e9ca2_result_delayed_u0=1'h0;
reg		reg_5874fe30_u0=1'h0;
reg		reg_3a9ed8da_u0=1'h0;
reg		reg_6f2cfbe7_result_delayed_result_delayed_u0=1'h0;
reg		reg_24a21cbf_result_delayed_result_delayed_u0=1'h0;
reg		reg_7ffc667d_result_delayed_result_delayed_u0=1'h0;
reg		reg_2efcd75c_result_delayed_u0=1'h0;
reg		reg_1796d9d9_u0=1'h0;
reg		reg_58a2a0e3_result_delayed_u0=1'h0;
reg		reg_04da25b8_result_delayed_u0=1'h0;
reg		reg_00246672_u0=1'h0;
reg		reg_6ec6926a_result_delayed_u0=1'h0;
reg		reg_32c8d37c_result_delayed_u0=1'h0;
reg		reg_0b8053fe_result_delayed_result_delayed_u0=1'h0;
reg		reg_0ee3ba53_result_delayed_result_delayed_u0=1'h0;
reg		reg_2976ab2a_u0=1'h0;
reg		reg_1fa5ca42_result_delayed_u0=1'h0;
reg		reg_1457ec7b_result_delayed_u0=1'h0;
reg		reg_68d00eb5_u0=1'h0;
reg		reg_68ca4866_result_delayed_u0=1'h0;
reg		reg_39c815b1_result_delayed_u0=1'h0;
reg		reg_1623704a_u0=1'h0;
reg		reg_5451da38_u0=1'h0;
reg		reg_7d510c70_result_delayed_u0=1'h0;
reg		reg_1036257e_result_delayed_u0=1'h0;
reg		reg_18e93e99_u0=1'h0;
reg		reg_7999bbe8_u0=1'h0;
reg		reg_1418995e_result_delayed_u0=1'h0;
reg		reg_677157b7_result_delayed_u0=1'h0;
reg		reg_4c7e6a09_u0=1'h0;
reg		reg_53090f63_result_delayed_u0=1'h0;
reg		reg_05b030d6_result_delayed_result_delayed_u0=1'h0;
reg		reg_4235f44a_u0=1'h0;
reg		reg_142b80f2_result_delayed_u0=1'h0;
reg		reg_09e28b61_u0=1'h0;
reg		reg_227958fa_u0=1'h0;
reg		reg_06efce9a_result_delayed_result_delayed_u0=1'h0;
reg		reg_52bc0089_result_delayed_u0=1'h0;
reg		reg_4e1c133b_result_delayed_result_delayed_u0=1'h0;
reg		reg_6028598b_result_delayed_result_delayed_u0=1'h0;
reg		reg_7bd0a7f4_result_delayed_u0=1'h0;
reg		reg_4d3893b7_u0=1'h0;
reg		reg_4235f44a_result_delayed_u0=1'h0;
reg		reg_690deb9c_u0=1'h0;
reg		reg_1ea77ba6_result_delayed_u0=1'h0;
reg		reg_1418995e_result_delayed_result_delayed_u0=1'h0;
reg		reg_18ff3a6a_u0=1'h0;
reg		reg_2ed4804d_u0=1'h0;
reg		reg_39c815b1_result_delayed_result_delayed_u0=1'h0;
reg		reg_640f5a91_u0=1'h0;
reg		reg_1ad50076_u0=1'h0;
reg		reg_1c1149c7_result_delayed_u0=1'h0;
reg		reg_4cc74cbd_result_delayed_result_delayed_u0=1'h0;
reg		reg_0f726638_result_delayed_u0=1'h0;
reg		reg_0a3ee092_u0=1'h0;
reg		reg_5451da38_result_delayed_u0=1'h0;
reg		reg_1fa5ca42_result_delayed_result_delayed_u0=1'h0;
reg		reg_4df0fb45_u0=1'h0;
reg		reg_6092b844_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_64049807_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_258244c0_result_delayed_u0=1'h0;
reg		reg_1457ec7b_result_delayed_result_delayed_u0=1'h0;
reg		reg_0b8053fe_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_1a0fb632_result_delayed_result_delayed_u0=1'h0;
reg		reg_3c2e9ca2_result_delayed_result_delayed_u0=1'h0;
reg		reg_0076a506_result_delayed_u0=1'h0;
reg		reg_75fb999e_result_delayed_u0=1'h0;
reg		reg_15c73839_result_delayed_u0=1'h0;
reg		reg_2f2401f0_u0=1'h0;
reg		reg_4235f44a_result_delayed_result_delayed_u0=1'h0;
reg		reg_576a3720_result_delayed_u0=1'h0;
reg		reg_7723f5fb_u0=1'h0;
reg		reg_426d8380_result_delayed_u0=1'h0;
reg		reg_26133792_result_delayed_u0=1'h0;
reg		reg_4d3893b7_result_delayed_u0=1'h0;
reg		reg_228ef2dc_result_delayed_u0=1'h0;
reg		reg_43da3530_u0=1'h0;
reg		reg_22603c8b_u0=1'h0;
reg		reg_21c538b9_result_delayed_u0=1'h0;
reg		reg_677157b7_result_delayed_result_delayed_u0=1'h0;
reg		reg_576a3720_result_delayed_result_delayed_u0=1'h0;
reg		reg_304f02b2_u0=1'h0;
reg		reg_0986382d_result_delayed_u0=1'h0;
reg		reg_6d17e172_result_delayed_u0=1'h0;
reg		reg_735b3058_u0=1'h0;
reg		reg_24a21cbf_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_201eb03b_result_delayed_u0=1'h0;
reg		reg_0bcf08c6_u0=1'h0;
reg		reg_747c90de_result_delayed_result_delayed_u0=1'h0;
reg		reg_0a6a1b0e_result_delayed_u0=1'h0;
reg		reg_2f9dd090_u0=1'h0;
reg		reg_30e8bfe6_u0=1'h0;
reg		reg_445ccdaa_result_delayed_u0=1'h0;
reg		reg_55edd085_result_delayed_u0=1'h0;
reg		reg_7807eb12_u0=1'h0;
reg		reg_1098e4cf_result_delayed_u0=1'h0;
reg		reg_242facb3_result_delayed_result_delayed_u0=1'h0;
reg		reg_77d7ef15_result_delayed_result_delayed_u0=1'h0;
reg		reg_7723f5fb_result_delayed_u0=1'h0;
reg		reg_0b769204_result_delayed_u0=1'h0;
reg		reg_367fcb5d_result_delayed_u0=1'h0;
reg		reg_387904fe_result_delayed_u0=1'h0;
reg		reg_104b8d92_result_delayed_u0=1'h0;
reg		reg_2537f8df_result_delayed_u0=1'h0;
reg		reg_04a57b8c_u0=1'h0;
reg		reg_2f9dd090_result_delayed_u0=1'h0;
reg		reg_7d61464a_u0=1'h0;
reg		reg_4235f44a_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_343e0093_result_delayed_u0=1'h0;
reg		reg_77668746_result_delayed_result_delayed_u0=1'h0;
reg		reg_00af20e1_result_delayed_u0=1'h0;
reg		reg_35c4a85b_result_delayed_u0=1'h0;
reg		reg_64daf8c4_result_delayed_u0=1'h0;
reg		reg_18ad0cb7_result_delayed_u0=1'h0;
reg		reg_68801c52_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_49242595_result_delayed_u0=1'h0;
reg		reg_1680ee34_result_delayed_u0=1'h0;
reg		reg_2c8dcfcc_u0=1'h0;
reg		reg_54ef10cf_result_delayed_u0=1'h0;
reg		reg_35d48481_result_delayed_u0=1'h0;
reg		reg_36ce22d8_result_delayed_u0=1'h0;
reg		reg_0425c0a1_result_delayed_u0=1'h0;
reg		reg_4a77e6f2_result_delayed_u0=1'h0;
reg		reg_5650d91a_u0=1'h0;
reg		reg_796241e6_result_delayed_u0=1'h0;
reg		reg_08eb52d0_result_delayed_u0=1'h0;
reg		reg_6a79fa17_result_delayed_u0=1'h0;
reg		reg_32a37dec_u0=1'h0;
reg		reg_38d95389_u0=1'h0;
reg		reg_70b8aa8a_result_delayed_u0=1'h0;
reg		reg_44a5d7f1_u0=1'h0;
reg		reg_5674bffb_result_delayed_u0=1'h0;
reg		reg_4769eae6_result_delayed_u0=1'h0;
reg		reg_4ffb5ab4_result_delayed_result_delayed_u0=1'h0;
reg		reg_441fe928_result_delayed_u0=1'h0;
wire		and_u2220_u0;
reg		reg_0a6a1b0e_result_delayed_result_delayed_u0=1'h0;
reg		reg_6bf613ee_result_delayed_u0=1'h0;
reg		reg_710efd1b_result_delayed_u0=1'h0;
reg		reg_1dd4f561_result_delayed_result_delayed_u0=1'h0;
reg		reg_09302a5b_u0=1'h0;
reg		reg_18e93e99_result_delayed_u0=1'h0;
wire		or_u690_u0;
wire		mux_u224;
reg		reg_0b8053fe_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_70b8aa8a_result_delayed_result_delayed_u0=1'h0;
reg		reg_227958fa_result_delayed_u0=1'h0;
reg		reg_382aec0c_result_delayed_result_delayed_u0=1'h0;
reg		reg_0fa7db18_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_09408e3d_u0=1'h0;
reg		reg_6092b844_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_4bbdc680_result_delayed_u0=1'h0;
reg		reg_13cde2f7_result_delayed_u0=1'h0;
reg		reg_343e0093_result_delayed_result_delayed_u0=1'h0;
reg		reg_7999bbe8_result_delayed_u0=1'h0;
reg		reg_4e289baa_result_delayed_u0=1'h0;
reg		reg_1a79d7d6_result_delayed_u0=1'h0;
reg		reg_1dd4f561_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_1a837eb0_result_delayed_u0=1'h0;
reg		reg_7bfae876_u0=1'h0;
reg		reg_7d46a529_result_delayed_u0=1'h0;
reg		reg_180dc380_u0=1'h0;
reg		reg_3a9ed8da_result_delayed_u0=1'h0;
reg		reg_70b8aa8a_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_32c8d37c_result_delayed_result_delayed_u0=1'h0;
reg		reg_64789d0a_result_delayed_u0=1'h0;
reg		reg_42536b9e_result_delayed_u0=1'h0;
reg		reg_229d1ee4_result_delayed_result_delayed_u0=1'h0;
reg		reg_1cd8b4df_result_delayed_u0=1'h0;
reg		reg_06dc9aa2_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_6f9e56f4_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_304f02b2_result_delayed_u0=1'h0;
reg		reg_5ee7823f_result_delayed_u0=1'h0;
reg		reg_6df7e814_result_delayed_result_delayed_u0=1'h0;
reg		reg_4a5adf10_result_delayed_result_delayed_u0=1'h0;
reg		reg_18ff3a6a_result_delayed_u0=1'h0;
reg		reg_4ffb5ab4_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_5e4d335d_result_delayed_result_delayed_u0=1'h0;
reg		reg_528f4535_u0=1'h0;
reg		reg_242facb3_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_00246672_result_delayed_u0=1'h0;
reg		reg_10810426_result_delayed_u0=1'h0;
reg		reg_09e28b61_result_delayed_u0=1'h0;
reg		reg_7a05baae_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_0f5456f1_result_delayed_u0=1'h0;
reg		reg_710f71fd_result_delayed_result_delayed_u0=1'h0;
reg		reg_426d8380_result_delayed_result_delayed_u0=1'h0;
reg		reg_6d759d56_result_delayed_result_delayed_u0=1'h0;
reg		reg_09e28b61_result_delayed_result_delayed_u0=1'h0;
reg		reg_640dac03_result_delayed_u0=1'h0;
reg		reg_2a321227_result_delayed_u0=1'h0;
reg		reg_2c8dcfcc_result_delayed_u0=1'h0;
reg		reg_6dec38b5_result_delayed_u0=1'h0;
reg		reg_5bc0cf31_result_delayed_result_delayed_u0=1'h0;
reg		reg_02369e1a_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_424e119f_u0=1'h0;
reg		reg_5c7b4c7d_result_delayed_result_delayed_u0=1'h0;
reg		reg_070292d1_result_delayed_u0=1'h0;
reg		reg_7e3e122c_result_delayed_u0=1'h0;
reg		reg_05b030d6_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_405c3132_result_delayed_u0=1'h0;
reg		reg_4a77e6f2_result_delayed_result_delayed_u0=1'h0;
reg		reg_0b38372d_result_delayed_result_delayed_u0=1'h0;
reg		reg_0d9b29cf_result_delayed_u0=1'h0;
reg		reg_5ee7823f_result_delayed_result_delayed_u0=1'h0;
reg		reg_2f9dd090_result_delayed_result_delayed_u0=1'h0;
reg		reg_1098e4cf_result_delayed_result_delayed_u0=1'h0;
reg		reg_39d6e99f_result_delayed_u0=1'h0;
reg		reg_7d231906_result_delayed_u0=1'h0;
reg		reg_47aed7f7_result_delayed_u0=1'h0;
reg		reg_104b8d92_result_delayed_result_delayed_u0=1'h0;
reg		reg_1dce6126_result_delayed_u0=1'h0;
reg		reg_183f91d8_result_delayed_u0=1'h0;
reg		reg_68e2082a_result_delayed_u0=1'h0;
reg		reg_64daf8c4_result_delayed_result_delayed_u0=1'h0;
reg		reg_76ad5fc6_result_delayed_u0=1'h0;
reg		reg_06efce9a_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_6dec38b5_result_delayed_result_delayed_u0=1'h0;
reg		reg_68ca4866_result_delayed_result_delayed_u0=1'h0;
reg		reg_2efcd75c_result_delayed_result_delayed_u0=1'h0;
reg		reg_6320b243_result_delayed_result_delayed_u0=1'h0;
reg		reg_2d8f78b3_result_delayed_u0=1'h0;
reg		reg_0f7cf45c_u0=1'h0;
wire		or_u691_u0;
wire	[31:0]	mux_u225_u0;
reg		reg_0f7cf45c_result_delayed_u0=1'h0;
wire		or_u692_u0;
wire		or_u693_u0;
wire		and_u2221_u0;
wire		or_u694_u0;
reg		reg_1f5cf7c4_u0=1'h0;
wire		and_u2222_u0;
reg		reg_1f5cf7c4_result_delayed_u0=1'h0;
reg		reg_0f7cf45c_result_delayed_result_delayed_u0=1'h0;
wire		or_u695_u0;
wire		mux_u226_u0;
wire		or_u696_u0;
wire		and_u2223_u0;
reg		reg_1769529a_u0=1'h0;
wire		or_u697_u0;
wire		and_u2224_u0;
wire		equals_u118;
wire signed	[31:0]	equals_u118_a_signed;
wire signed	[31:0]	equals_u118_b_signed;
wire		and_u2225_u0;
wire		and_u2226_u0;
wire		not_u409_u0;
wire		not_u410_u0;
wire		and_u2227_u0;
wire		and_u2228_u0;
wire		lessThan_u51;
wire signed	[31:0]	lessThan_u51_b_signed;
wire signed	[31:0]	lessThan_u51_a_signed;
wire		not_u411_u0;
wire		and_u2229_u0;
wire		and_u2230_u0;
wire		and_u2231_u0;
wire		not_u412_u0;
wire		and_u2232_u0;
wire	[31:0]	add;
wire		and_u2233_u0;
wire		simplePinWrite_u368;
wire	[15:0]	simplePinWrite_u369;
wire	[15:0]	simplePinWrite_u370;
wire	[31:0]	add_u167;
reg	[15:0]	syncEnable_u317=16'h0;
wire	[15:0]	mux_u227_u0;
reg		reg_3543084e_u0=1'h0;
wire		and_u2234_u0;
reg		and_delayed_u145=1'h0;
reg	[15:0]	syncEnable_u318_u0=16'h0;
wire		and_u2235_u0;
reg	[31:0]	syncEnable_u319_u0=32'h0;
reg	[15:0]	syncEnable_u320_u0=16'h0;
wire	[15:0]	mux_u228_u0;
reg		reg_394c9807_u0=1'h0;
wire	[31:0]	mux_u229_u0;
wire		and_u2236_u0;
reg		reg_5a8744bc_u0=1'h0;
wire		and_u2237_u0;
wire	[31:0]	mux_u230_u0;
reg		reg_371d79bc_u0=1'h0;
wire		and_u2238_u0;
reg	[31:0]	syncEnable_u321_u0=32'h0;
wire		and_u2239_u0;
reg	[15:0]	syncEnable_u322_u0=16'h0;
reg		and_delayed_u146_u0=1'h0;
wire	[15:0]	mux_u231_u0;
wire	[31:0]	mux_u232_u0;
wire		and_u2240_u0;
wire		and_u2241_u0;
wire	[15:0]	mux_u233_u0;
reg		and_delayed_u147_u0=1'h0;
reg	[15:0]	syncEnable_u323_u0=16'h0;
reg		and_delayed_u148_u0=1'h0;
reg	[31:0]	syncEnable_u324_u0=32'h0;
wire	[31:0]	mux_u234_u0;
wire		or_u698_u0;
wire		or_u699_u0;
wire		mux_u235_u0;
wire		mux_u236_u0;
wire		or_u700_u0;
reg		block_GO_delayed_u8=1'h0;
reg	[15:0]	latch_2c039393_reg=16'h0;
wire	[15:0]	latch_2c039393_out;
reg	[31:0]	latch_36791ce1_reg=32'h0;
wire	[31:0]	latch_36791ce1_out;
wire	[31:0]	mux_u237_u0;
wire		or_u701_u0;
wire		and_u2242_u0;
reg	[15:0]	fbReg_Out1Portvalue_u1=16'h0;
reg		syncEnable_u325_u0=1'h0;
wire	[15:0]	mux_u238_u0;
wire		or_u702_u0;
reg	[31:0]	fbReg_temp_fsmOldState_resized_HH2_xy_4_u0=32'h0;
wire	[31:0]	mux_u239_u0;
reg		loopControl_u5=1'h0;
wire		or_u703_u0;
wire		or_u704_u0;
wire		mux_u240_u0;
reg		reg_01da6964_u0=1'h0;
wire		or_u705_u0;
wire		mux_u241_u0;
wire		or_u706_u0;
wire	[31:0]	mux_u242_u0;
wire		or_u707_u0;
wire	[31:0]	mux_u243_u0;
reg		reg_1c62611c_u0=1'h0;
assign lessThan_a_unsigned=port_038b3c60_;
assign lessThan_b_unsigned=16'h80;
assign lessThan=lessThan_a_unsigned<lessThan_b_unsigned;
assign equals_a_unsigned=port_038b3c60_;
assign equals_b_unsigned=16'h80;
assign equals=equals_a_unsigned==equals_b_unsigned;
assign lessThan_u50_a_unsigned=port_7451eb09_;
assign lessThan_u50_b_unsigned=16'h4;
assign lessThan_u50=lessThan_u50_a_unsigned<lessThan_u50_b_unsigned;
assign andOp=equals&lessThan_u50;
assign equals_u116_a_unsigned=port_7451eb09_;
assign equals_u116_b_unsigned=16'h4;
assign equals_u116=equals_u116_a_unsigned==equals_u116_b_unsigned;
assign equals_u117_a_signed={31'b0, port_768be70f_};
assign equals_u117_b_signed=32'h0;
assign equals_u117=equals_u117_a_signed==equals_u117_b_signed;
assign and_u2210_u0=and_u2242_u0&not_u405_u0;
assign not_u405_u0=~equals_u117;
assign and_u2211_u0=and_u2242_u0&equals_u117;
assign andOp_u133=lessThan&port_1bbb1093_;
assign not_u406_u0=~andOp_u133;
assign and_u2212_u0=and_u2223_u0&not_u406_u0;
assign and_u2213_u0=and_u2223_u0&andOp_u133;
assign simplePinWrite=and_u2221_u0&{1{and_u2221_u0}};
assign not_u407_u0=~andOp;
assign and_u2214_u0=and_u2222_u0&andOp;
assign and_u2215_u0=and_u2222_u0&not_u407_u0;
assign simplePinWrite_u366=and_u2220_u0&{1{and_u2220_u0}};
assign and_u2216_u0=and_u2219_u0&equals_u116;
assign not_u408_u0=~equals_u116;
assign and_u2217_u0=and_u2219_u0&not_u408_u0;
assign simplePinWrite_u367=and_u2218_u0&{1{and_u2218_u0}};
assign and_u2218_u0=and_u2216_u0&and_u2219_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_62bcd2be_u0<=1'h0;
else reg_62bcd2be_u0<=reg_31a64119_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_64049807_u0<=1'h0;
else reg_64049807_u0<=reg_0ee3ba53_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5c7b4c7d_u0<=1'h0;
else reg_5c7b4c7d_u0<=reg_228ef2dc_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1cd8b4df_u0<=1'h0;
else reg_1cd8b4df_u0<=reg_30e4f8f8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_640dac03_u0<=1'h0;
else reg_640dac03_u0<=reg_7d61464a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7e3e122c_u0<=1'h0;
else reg_7e3e122c_u0<=reg_38645974_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0b38372d_u0<=1'h0;
else reg_0b38372d_u0<=reg_532c937d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_710efd1b_u0<=1'h0;
else reg_710efd1b_u0<=reg_43da3530_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2a321227_u0<=1'h0;
else reg_2a321227_u0<=reg_183f91d8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_36ce22d8_u0<=1'h0;
else reg_36ce22d8_u0<=reg_66565274_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6bf613ee_u0<=1'h0;
else reg_6bf613ee_u0<=reg_4c9f1046_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_18ad0cb7_u0<=1'h0;
else reg_18ad0cb7_u0<=reg_34d4a805_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_30e4f8f8_u0<=1'h0;
else reg_30e4f8f8_u0<=reg_5e188306_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_24a21cbf_u0<=1'h0;
else reg_24a21cbf_u0<=reg_1f1eb78a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_64daf8c4_u0<=1'h0;
else reg_64daf8c4_u0<=reg_09a32d61_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_54ef10cf_u0<=1'h0;
else reg_54ef10cf_u0<=reg_2c1074d0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_77668746_u0<=1'h0;
else reg_77668746_u0<=reg_337b1691_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_77668746_result_delayed_u0<=1'h0;
else reg_77668746_result_delayed_u0<=reg_77668746_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_66565274_u0<=1'h0;
else reg_66565274_u0<=reg_0320d63a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6d759d56_u0<=1'h0;
else reg_6d759d56_u0<=reg_528f4535_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7bd0a7f4_u0<=1'h0;
else reg_7bd0a7f4_u0<=reg_6d17e172_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_201eb03b_u0<=1'h0;
else reg_201eb03b_u0<=reg_027e723d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7d231906_u0<=1'h0;
else reg_7d231906_u0<=reg_1ad50076_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_42b58a90_u0<=1'h0;
else reg_42b58a90_u0<=reg_5101c4c6_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_382aec0c_u0<=1'h0;
else reg_382aec0c_u0<=reg_4cc74cbd_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1457ec7b_u0<=1'h0;
else reg_1457ec7b_u0<=reg_06efce9a_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_02369e1a_u0<=1'h0;
else reg_02369e1a_u0<=reg_42b58a90_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6848807a_u0<=1'h0;
else reg_6848807a_u0<=reg_66c4e649_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1a837eb0_u0<=1'h0;
else reg_1a837eb0_u0<=reg_677157b7_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_45a11597_u0<=1'h0;
else reg_45a11597_u0<=reg_2a60e877_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_774ab77d_u0<=1'h0;
else reg_774ab77d_u0<=reg_7a05baae_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_62921ea8_u0<=1'h0;
else reg_62921ea8_u0<=reg_2f2401f0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0034740f_u0<=1'h0;
else reg_0034740f_u0<=reg_579a33fd_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1a0fb632_u0<=1'h0;
else reg_1a0fb632_u0<=reg_03b6ff07_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_061a1224_u0<=1'h0;
else reg_061a1224_u0<=reg_6320b243_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_58a2a0e3_u0<=1'h0;
else reg_58a2a0e3_u0<=reg_44a5d7f1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_027e723d_u0<=1'h0;
else reg_027e723d_u0<=reg_5c7b4c7d_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_39d6e99f_u0<=1'h0;
else reg_39d6e99f_u0<=reg_650388ee_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_576a3720_u0<=1'h0;
else reg_576a3720_u0<=reg_18e93e99_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_30e4f8f8_result_delayed_u0<=1'h0;
else reg_30e4f8f8_result_delayed_u0<=reg_30e4f8f8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00af20e1_u0<=1'h0;
else reg_00af20e1_u0<=reg_774ab77d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_532c937d_u0<=1'h0;
else reg_532c937d_u0<=reg_5ee7823f_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_228ef2dc_u0<=1'h0;
else reg_228ef2dc_u0<=reg_3c2e9ca2_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_02369e1a_result_delayed_u0<=1'h0;
else reg_02369e1a_result_delayed_u0<=reg_02369e1a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0d9b29cf_u0<=1'h0;
else reg_0d9b29cf_u0<=reg_6ec6926a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1098e4cf_u0<=1'h0;
else reg_1098e4cf_u0<=reg_5046f020_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_47aed7f7_u0<=1'h0;
else reg_47aed7f7_u0<=reg_0986382d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0ced50b0_u0<=1'h0;
else reg_0ced50b0_u0<=reg_09069cf0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6d17e172_u0<=1'h0;
else reg_6d17e172_u0<=reg_1dff8122_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_75fb999e_u0<=1'h0;
else reg_75fb999e_u0<=reg_42536b9e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5046f020_u0<=1'h0;
else reg_5046f020_u0<=reg_48ad5013_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_579a33fd_u0<=1'h0;
else reg_579a33fd_u0<=reg_1036257e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_53090f63_u0<=1'h0;
else reg_53090f63_u0<=reg_62b86a49_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_38a628ca_u0<=1'h0;
else reg_38a628ca_u0<=reg_010c659c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6a79fa17_u0<=1'h0;
else reg_6a79fa17_u0<=reg_64e0b984_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_02369e1a_result_delayed_result_delayed_u0<=1'h0;
else reg_02369e1a_result_delayed_result_delayed_u0<=reg_02369e1a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7d46a529_u0<=1'h0;
else reg_7d46a529_u0<=reg_09e28b61_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_06efce9a_u0<=1'h0;
else reg_06efce9a_u0<=reg_15c73839_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1a0fb632_result_delayed_u0<=1'h0;
else reg_1a0fb632_result_delayed_u0<=reg_1a0fb632_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_24a21cbf_result_delayed_u0<=1'h0;
else reg_24a21cbf_result_delayed_u0<=reg_24a21cbf_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4cd00ca8_u0<=1'h0;
else reg_4cd00ca8_u0<=reg_10810426_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_39c815b1_u0<=1'h0;
else reg_39c815b1_u0<=reg_227958fa_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_229d1ee4_u0<=1'h0;
else reg_229d1ee4_u0<=reg_22603c8b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4cc74cbd_u0<=1'h0;
else reg_4cc74cbd_u0<=reg_0f2ec27d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6d923de9_u0<=1'h0;
else reg_6d923de9_u0<=and_u2219_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0b8053fe_u0<=1'h0;
else reg_0b8053fe_u0<=reg_7bfae876_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_06dc9aa2_u0<=1'h0;
else reg_06dc9aa2_u0<=reg_35da3503_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_796241e6_u0<=1'h0;
else reg_796241e6_u0<=reg_2add40ec_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0425c0a1_u0<=1'h0;
else reg_0425c0a1_u0<=reg_30e8bfe6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4a77e6f2_u0<=1'h0;
else reg_4a77e6f2_u0<=reg_0076a506_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_387904fe_u0<=1'h0;
else reg_387904fe_u0<=reg_02369e1a_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3c2e9ca2_u0<=1'h0;
else reg_3c2e9ca2_u0<=reg_0b8053fe_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_66c4e649_u0<=1'h0;
else reg_66c4e649_u0<=reg_13b25f04_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_010c659c_u0<=1'h0;
else reg_010c659c_u0<=reg_1623704a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_774ab77d_result_delayed_u0<=1'h0;
else reg_774ab77d_result_delayed_u0<=reg_774ab77d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4cc74cbd_result_delayed_u0<=1'h0;
else reg_4cc74cbd_result_delayed_u0<=reg_4cc74cbd_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1f1eb78a_u0<=1'h0;
else reg_1f1eb78a_u0<=reg_7010ad01_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0346d3d3_u0<=1'h0;
else reg_0346d3d3_u0<=reg_0a6a1b0e_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6a895611_u0<=1'h0;
else reg_6a895611_u0<=reg_18ad0cb7_result_delayed_u0;
end
assign and_u2219_u0=and_u2215_u0&and_u2222_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_242facb3_u0<=1'h0;
else reg_242facb3_u0<=reg_439b9ebb_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_747c90de_u0<=1'h0;
else reg_747c90de_u0<=reg_4ca109c7_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_38a0bc03_u0<=1'h0;
else reg_38a0bc03_u0<=reg_29ad1d65_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_31615dc2_u0<=1'h0;
else reg_31615dc2_u0<=reg_2d8f78b3_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_10810426_u0<=1'h0;
else reg_10810426_u0<=reg_7e3e122c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a05baae_u0<=1'h0;
else reg_7a05baae_u0<=reg_75ddf3cd_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_68ca4866_u0<=1'h0;
else reg_68ca4866_u0<=reg_1ea77ba6_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6ec6926a_u0<=1'h0;
else reg_6ec6926a_u0<=reg_1796d9d9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_343e0093_u0<=1'h0;
else reg_343e0093_u0<=reg_5e4d335d_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0b8053fe_result_delayed_u0<=1'h0;
else reg_0b8053fe_result_delayed_u0<=reg_0b8053fe_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0ee3ba53_u0<=1'h0;
else reg_0ee3ba53_u0<=reg_2ea3b7cc_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2894b025_u0<=1'h0;
else reg_2894b025_u0<=reg_56b4ebc1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_03b6ff07_u0<=1'h0;
else reg_03b6ff07_u0<=reg_7723f5fb_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_49242595_u0<=1'h0;
else reg_49242595_u0<=reg_24a21cbf_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1680ee34_u0<=1'h0;
else reg_1680ee34_u0<=reg_14de3123_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1dd4f561_u0<=1'h0;
else reg_1dd4f561_u0<=reg_01a00b9a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_13b25f04_u0<=1'h0;
else reg_13b25f04_u0<=reg_22f13343_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_06efce9a_result_delayed_u0<=1'h0;
else reg_06efce9a_result_delayed_u0<=reg_06efce9a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_48ad5013_u0<=1'h0;
else reg_48ad5013_u0<=reg_6848807a_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1c7bd8c5_u0<=1'h0;
else reg_1c7bd8c5_u0<=reg_62921ea8_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_31a64119_u0<=1'h0;
else reg_31a64119_u0<=reg_5874fe30_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0fa7db18_u0<=1'h0;
else reg_0fa7db18_u0<=reg_29984143_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2c1074d0_u0<=1'h0;
else reg_2c1074d0_u0<=reg_1a837eb0_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_09a32d61_u0<=1'h0;
else reg_09a32d61_u0<=reg_04da25b8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_77d7ef15_u0<=1'h0;
else reg_77d7ef15_u0<=reg_3a15fb72_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_677157b7_u0<=1'h0;
else reg_677157b7_u0<=reg_0ced50b0_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_68e2082a_u0<=1'h0;
else reg_68e2082a_u0<=reg_4a3f86cf_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_29ad1d65_u0<=1'h0;
else reg_29ad1d65_u0<=reg_4a5adf10_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6f2cfbe7_u0<=1'h0;
else reg_6f2cfbe7_u0<=reg_7ffc667d_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_34d4a805_u0<=1'h0;
else reg_34d4a805_u0<=reg_061a1224_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_68801c52_u0<=1'h0;
else reg_68801c52_u0<=reg_0530331a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6092b844_u0<=1'h0;
else reg_6092b844_u0<=reg_6c7e010b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5ee7823f_u0<=1'h0;
else reg_5ee7823f_u0<=reg_1680ee34_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6d759d56_result_delayed_u0<=1'h0;
else reg_6d759d56_result_delayed_u0<=reg_6d759d56_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_35da3503_u0<=1'h0;
else reg_35da3503_u0<=reg_6a895611_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4c9f1046_u0<=1'h0;
else reg_4c9f1046_u0<=reg_258244c0_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_142b80f2_u0<=1'h0;
else reg_142b80f2_u0<=reg_24232921_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_29984143_u0<=1'h0;
else reg_29984143_u0<=reg_33b2aabd_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1dff8122_u0<=1'h0;
else reg_1dff8122_u0<=reg_40fef52d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_229d1ee4_result_delayed_u0<=1'h0;
else reg_229d1ee4_result_delayed_u0<=reg_229d1ee4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1dce6126_u0<=1'h0;
else reg_1dce6126_u0<=reg_09302a5b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6848807a_result_delayed_u0<=1'h0;
else reg_6848807a_result_delayed_u0<=reg_6848807a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_42b58a90_result_delayed_u0<=1'h0;
else reg_42b58a90_result_delayed_u0<=reg_42b58a90_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4a3f86cf_u0<=1'h0;
else reg_4a3f86cf_u0<=reg_0346d3d3_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5a7e368e_u0<=1'h0;
else reg_5a7e368e_u0<=reg_6028598b_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_62921ea8_result_delayed_u0<=1'h0;
else reg_62921ea8_result_delayed_u0<=reg_62921ea8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5bc0cf31_u0<=1'h0;
else reg_5bc0cf31_u0<=reg_38a628ca_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6a895611_result_delayed_u0<=1'h0;
else reg_6a895611_result_delayed_u0<=reg_6a895611_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_62b86a49_u0<=1'h0;
else reg_62b86a49_u0<=reg_3f8e0a19_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4589457b_u0<=1'h0;
else reg_4589457b_u0<=reg_0034740f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_710f71fd_u0<=1'h0;
else reg_710f71fd_u0<=reg_0fa7db18_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6092b844_result_delayed_u0<=1'h0;
else reg_6092b844_result_delayed_u0<=reg_6092b844_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6f2cfbe7_result_delayed_u0<=1'h0;
else reg_6f2cfbe7_result_delayed_u0<=reg_6f2cfbe7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1ea77ba6_u0<=1'h0;
else reg_1ea77ba6_u0<=reg_62bcd2be_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_62921ea8_result_delayed_result_delayed_u0<=1'h0;
else reg_62921ea8_result_delayed_result_delayed_u0<=reg_62921ea8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_24232921_u0<=1'h0;
else reg_24232921_u0<=reg_28e37146_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_06dc9aa2_result_delayed_u0<=1'h0;
else reg_06dc9aa2_result_delayed_u0<=reg_06dc9aa2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_33b2aabd_u0<=1'h0;
else reg_33b2aabd_u0<=reg_0425c0a1_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5e4d335d_u0<=1'h0;
else reg_5e4d335d_u0<=reg_45a11597_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_38645974_u0<=1'h0;
else reg_38645974_u0<=reg_4589457b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7010ad01_u0<=1'h0;
else reg_7010ad01_u0<=reg_1dce6126_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0320d63a_u0<=1'h0;
else reg_0320d63a_u0<=reg_1cd8b4df_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5e188306_u0<=1'h0;
else reg_5e188306_u0<=reg_640dac03_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0fa7db18_result_delayed_u0<=1'h0;
else reg_0fa7db18_result_delayed_u0<=reg_0fa7db18_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_439b9ebb_u0<=1'h0;
else reg_439b9ebb_u0<=reg_4ec55fe6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7d510c70_u0<=1'h0;
else reg_7d510c70_u0<=reg_5451da38_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_367fcb5d_u0<=1'h0;
else reg_367fcb5d_u0<=reg_2894b025_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4ec55fe6_u0<=1'h0;
else reg_4ec55fe6_u0<=reg_0bcf08c6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0ced50b0_result_delayed_u0<=1'h0;
else reg_0ced50b0_result_delayed_u0<=reg_0ced50b0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4e1c133b_u0<=1'h0;
else reg_4e1c133b_u0<=reg_6092b844_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_061a1224_result_delayed_u0<=1'h0;
else reg_061a1224_result_delayed_u0<=reg_061a1224_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6092b844_result_delayed_result_delayed_u0<=1'h0;
else reg_6092b844_result_delayed_result_delayed_u0<=reg_6092b844_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_441fe928_u0<=1'h0;
else reg_441fe928_u0<=reg_35c4a85b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_13cde2f7_u0<=1'h0;
else reg_13cde2f7_u0<=reg_4cd00ca8_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2d8f78b3_u0<=1'h0;
else reg_2d8f78b3_u0<=reg_7d212c9a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4bbdc680_u0<=1'h0;
else reg_4bbdc680_u0<=reg_2976ab2a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_258244c0_u0<=1'h0;
else reg_258244c0_u0<=reg_104b8d92_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_06dc9aa2_result_delayed_result_delayed_u0<=1'h0;
else reg_06dc9aa2_result_delayed_result_delayed_u0<=reg_06dc9aa2_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_38a0bc03_result_delayed_u0<=1'h0;
else reg_38a0bc03_result_delayed_u0<=reg_38a0bc03_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1418995e_u0<=1'h0;
else reg_1418995e_u0<=reg_242facb3_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1036257e_u0<=1'h0;
else reg_1036257e_u0<=reg_2537f8df_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5e4d335d_result_delayed_u0<=1'h0;
else reg_5e4d335d_result_delayed_u0<=reg_5e4d335d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4a5adf10_u0<=1'h0;
else reg_4a5adf10_u0<=reg_150760de_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0f726638_u0<=1'h0;
else reg_0f726638_u0<=reg_1c1149c7_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4ffb5ab4_u0<=1'h0;
else reg_4ffb5ab4_u0<=reg_58a2a0e3_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6848807a_result_delayed_result_delayed_u0<=1'h0;
else reg_6848807a_result_delayed_result_delayed_u0<=reg_6848807a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0f2ec27d_u0<=1'h0;
else reg_0f2ec27d_u0<=reg_304f02b2_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_35d48481_u0<=1'h0;
else reg_35d48481_u0<=reg_1457ec7b_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6dec38b5_u0<=1'h0;
else reg_6dec38b5_u0<=reg_735b3058_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5bc0cf31_result_delayed_u0<=1'h0;
else reg_5bc0cf31_result_delayed_u0<=reg_5bc0cf31_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_64049807_result_delayed_u0<=1'h0;
else reg_64049807_result_delayed_u0<=reg_64049807_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_04da25b8_u0<=1'h0;
else reg_04da25b8_u0<=reg_2ed4804d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6320b243_u0<=1'h0;
else reg_6320b243_u0<=reg_0cc8a5bf_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0a6a1b0e_u0<=1'h0;
else reg_0a6a1b0e_u0<=and_u2220_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_747c90de_result_delayed_u0<=1'h0;
else reg_747c90de_result_delayed_u0<=reg_747c90de_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_64e0b984_u0<=1'h0;
else reg_64e0b984_u0<=reg_38a0bc03_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_42b58a90_result_delayed_result_delayed_u0<=1'h0;
else reg_42b58a90_result_delayed_result_delayed_u0<=reg_42b58a90_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_05b030d6_u0<=1'h0;
else reg_05b030d6_u0<=reg_53090f63_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4ca109c7_u0<=1'h0;
else reg_4ca109c7_u0<=reg_1a0fb632_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3a15fb72_u0<=1'h0;
else reg_3a15fb72_u0<=reg_5a7e368e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_55edd085_u0<=1'h0;
else reg_55edd085_u0<=reg_47aed7f7_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0034740f_result_delayed_u0<=1'h0;
else reg_0034740f_result_delayed_u0<=reg_0034740f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6f9e56f4_u0<=1'h0;
else reg_6f9e56f4_u0<=reg_76f5e34d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_76ad5fc6_u0<=1'h0;
else reg_76ad5fc6_u0<=reg_3ecadb64_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6320b243_result_delayed_u0<=1'h0;
else reg_6320b243_result_delayed_u0<=reg_6320b243_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1dd4f561_result_delayed_u0<=1'h0;
else reg_1dd4f561_result_delayed_u0<=reg_1dd4f561_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0b38372d_result_delayed_u0<=1'h0;
else reg_0b38372d_result_delayed_u0<=reg_0b38372d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_405c3132_u0<=1'h0;
else reg_405c3132_u0<=reg_382aec0c_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2ea3b7cc_u0<=1'h0;
else reg_2ea3b7cc_u0<=reg_2f9dd090_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0076a506_u0<=1'h0;
else reg_0076a506_u0<=reg_576a3720_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4a5adf10_result_delayed_u0<=1'h0;
else reg_4a5adf10_result_delayed_u0<=reg_4a5adf10_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0b769204_u0<=1'h0;
else reg_0b769204_u0<=reg_4e289baa_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_64789d0a_u0<=1'h0;
else reg_64789d0a_u0<=reg_51172316_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_56b4ebc1_u0<=1'h0;
else reg_56b4ebc1_u0<=reg_64049807_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6c7e010b_u0<=1'h0;
else reg_6c7e010b_u0<=reg_77d7ef15_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4ca109c7_result_delayed_u0<=1'h0;
else reg_4ca109c7_result_delayed_u0<=reg_4ca109c7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0cc8a5bf_u0<=1'h0;
else reg_0cc8a5bf_u0<=reg_222ee43c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_35da3503_result_delayed_u0<=1'h0;
else reg_35da3503_result_delayed_u0<=reg_35da3503_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_21c538b9_u0<=1'h0;
else reg_21c538b9_u0<=reg_08eb52d0_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6f9e56f4_result_delayed_u0<=1'h0;
else reg_6f9e56f4_result_delayed_u0<=reg_6f9e56f4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7ffc667d_u0<=1'h0;
else reg_7ffc667d_u0<=reg_7338c2c5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_26133792_u0<=1'h0;
else reg_26133792_u0<=reg_1418995e_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4e289baa_u0<=1'h0;
else reg_4e289baa_u0<=reg_32a37dec_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_579a33fd_result_delayed_u0<=1'h0;
else reg_579a33fd_result_delayed_u0<=reg_579a33fd_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_710f71fd_result_delayed_u0<=1'h0;
else reg_710f71fd_result_delayed_u0<=reg_710f71fd_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4cd00ca8_result_delayed_u0<=1'h0;
else reg_4cd00ca8_result_delayed_u0<=reg_4cd00ca8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_382aec0c_result_delayed_u0<=1'h0;
else reg_382aec0c_result_delayed_u0<=reg_382aec0c_u0;
end
assign or_u689_u0=reg_31615dc2_u0|reg_6d923de9_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_38a0bc03_result_delayed_result_delayed_u0<=1'h0;
else reg_38a0bc03_result_delayed_result_delayed_u0<=reg_38a0bc03_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4e1c133b_result_delayed_u0<=1'h0;
else reg_4e1c133b_result_delayed_u0<=reg_4e1c133b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5674bffb_u0<=1'h0;
else reg_5674bffb_u0<=reg_0f5456f1_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4769eae6_u0<=1'h0;
else reg_4769eae6_u0<=reg_387904fe_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a05baae_result_delayed_u0<=1'h0;
else reg_7a05baae_result_delayed_u0<=reg_7a05baae_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3f8e0a19_u0<=1'h0;
else reg_3f8e0a19_u0<=reg_7d510c70_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5c7b4c7d_result_delayed_u0<=1'h0;
else reg_5c7b4c7d_result_delayed_u0<=reg_5c7b4c7d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_45a11597_result_delayed_u0<=1'h0;
else reg_45a11597_result_delayed_u0<=reg_45a11597_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6c7e010b_result_delayed_u0<=1'h0;
else reg_6c7e010b_result_delayed_u0<=reg_6c7e010b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_242facb3_result_delayed_u0<=1'h0;
else reg_242facb3_result_delayed_u0<=reg_242facb3_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_35c4a85b_u0<=1'h0;
else reg_35c4a85b_u0<=reg_38d95389_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2efcd75c_u0<=1'h0;
else reg_2efcd75c_u0<=reg_35d48481_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_29984143_result_delayed_u0<=1'h0;
else reg_29984143_result_delayed_u0<=reg_29984143_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6028598b_u0<=1'h0;
else reg_6028598b_u0<=reg_7d46a529_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0f5456f1_u0<=1'h0;
else reg_0f5456f1_u0<=reg_2efcd75c_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_28e37146_u0<=1'h0;
else reg_28e37146_u0<=reg_424e119f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_42b58a90_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_42b58a90_result_delayed_result_delayed_result_delayed_u0<=reg_42b58a90_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_77d7ef15_result_delayed_u0<=1'h0;
else reg_77d7ef15_result_delayed_u0<=reg_77d7ef15_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4cd00ca8_result_delayed_result_delayed_u0<=1'h0;
else reg_4cd00ca8_result_delayed_result_delayed_u0<=reg_4cd00ca8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0986382d_u0<=1'h0;
else reg_0986382d_u0<=reg_64789d0a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3ecadb64_u0<=1'h0;
else reg_3ecadb64_u0<=reg_70b8aa8a_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1a79d7d6_u0<=1'h0;
else reg_1a79d7d6_u0<=reg_09408e3d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_22f13343_u0<=1'h0;
else reg_22f13343_u0<=reg_4e1c133b_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_32c8d37c_u0<=1'h0;
else reg_32c8d37c_u0<=reg_3a9ed8da_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4f367a8e_u0<=1'h0;
else reg_4f367a8e_u0<=reg_75fb999e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_76f5e34d_u0<=1'h0;
else reg_76f5e34d_u0<=reg_21c538b9_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0346d3d3_result_delayed_u0<=1'h0;
else reg_0346d3d3_result_delayed_u0<=reg_0346d3d3_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7d212c9a_u0<=1'h0;
else reg_7d212c9a_u0<=reg_195de36c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_64049807_result_delayed_result_delayed_u0<=1'h0;
else reg_64049807_result_delayed_result_delayed_u0<=reg_64049807_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5101c4c6_u0<=1'h0;
else reg_5101c4c6_u0<=reg_18ff3a6a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4589457b_result_delayed_u0<=1'h0;
else reg_4589457b_result_delayed_u0<=reg_4589457b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_02369e1a_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_02369e1a_result_delayed_result_delayed_result_delayed_u0<=reg_02369e1a_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a05baae_result_delayed_result_delayed_u0<=1'h0;
else reg_7a05baae_result_delayed_result_delayed_u0<=reg_7a05baae_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_42536b9e_u0<=1'h0;
else reg_42536b9e_u0<=reg_4d3893b7_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7010ad01_result_delayed_u0<=1'h0;
else reg_7010ad01_result_delayed_u0<=reg_7010ad01_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_40fef52d_u0<=1'h0;
else reg_40fef52d_u0<=reg_0b38372d_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_070292d1_u0<=1'h0;
else reg_070292d1_u0<=reg_0d9b29cf_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_42b58a90_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_42b58a90_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_42b58a90_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1c1149c7_u0<=1'h0;
else reg_1c1149c7_u0<=reg_1fbac5be_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6028598b_result_delayed_u0<=1'h0;
else reg_6028598b_result_delayed_u0<=reg_6028598b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_64049807_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_64049807_result_delayed_result_delayed_result_delayed_u0<=reg_64049807_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_150760de_u0<=1'h0;
else reg_150760de_u0<=reg_690deb9c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_104b8d92_u0<=1'h0;
else reg_104b8d92_u0<=reg_1c7bd8c5_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0ee3ba53_result_delayed_u0<=1'h0;
else reg_0ee3ba53_result_delayed_u0<=reg_0ee3ba53_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7ffc667d_result_delayed_u0<=1'h0;
else reg_7ffc667d_result_delayed_u0<=reg_7ffc667d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_38a628ca_result_delayed_u0<=1'h0;
else reg_38a628ca_result_delayed_u0<=reg_38a628ca_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6df7e814_u0<=1'h0;
else reg_6df7e814_u0<=reg_1a79d7d6_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5101c4c6_result_delayed_u0<=1'h0;
else reg_5101c4c6_result_delayed_u0<=reg_5101c4c6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1fa5ca42_u0<=1'h0;
else reg_1fa5ca42_u0<=reg_5df79fda_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_183f91d8_u0<=1'h0;
else reg_183f91d8_u0<=reg_142b80f2_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2537f8df_u0<=1'h0;
else reg_2537f8df_u0<=reg_68d00eb5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_337b1691_u0<=1'h0;
else reg_337b1691_u0<=reg_4bbdc680_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_426d8380_u0<=1'h0;
else reg_426d8380_u0<=reg_0a3ee092_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_650388ee_u0<=1'h0;
else reg_650388ee_u0<=reg_55edd085_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2894b025_result_delayed_u0<=1'h0;
else reg_2894b025_result_delayed_u0<=reg_2894b025_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_48ad5013_result_delayed_u0<=1'h0;
else reg_48ad5013_result_delayed_u0<=reg_48ad5013_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_68801c52_result_delayed_u0<=1'h0;
else reg_68801c52_result_delayed_u0<=reg_68801c52_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_09069cf0_u0<=1'h0;
else reg_09069cf0_u0<=reg_4a77e6f2_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_445ccdaa_u0<=1'h0;
else reg_445ccdaa_u0<=reg_6d759d56_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_14de3123_u0<=1'h0;
else reg_14de3123_u0<=reg_54ef10cf_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_62bcd2be_result_delayed_u0<=1'h0;
else reg_62bcd2be_result_delayed_u0<=reg_62bcd2be_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7338c2c5_u0<=1'h0;
else reg_7338c2c5_u0<=reg_796241e6_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_15c73839_u0<=1'h0;
else reg_15c73839_u0<=reg_4f367a8e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_51172316_u0<=1'h0;
else reg_51172316_u0<=reg_49242595_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1fbac5be_u0<=1'h0;
else reg_1fbac5be_u0<=reg_13cde2f7_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4ffb5ab4_result_delayed_u0<=1'h0;
else reg_4ffb5ab4_result_delayed_u0<=reg_4ffb5ab4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5a7e368e_result_delayed_u0<=1'h0;
else reg_5a7e368e_result_delayed_u0<=reg_5a7e368e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_38a628ca_result_delayed_result_delayed_u0<=1'h0;
else reg_38a628ca_result_delayed_result_delayed_u0<=reg_38a628ca_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6f9e56f4_result_delayed_result_delayed_u0<=1'h0;
else reg_6f9e56f4_result_delayed_result_delayed_u0<=reg_6f9e56f4_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_75ddf3cd_u0<=1'h0;
else reg_75ddf3cd_u0<=reg_06dc9aa2_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_222ee43c_u0<=1'h0;
else reg_222ee43c_u0<=reg_6f2cfbe7_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_24232921_result_delayed_u0<=1'h0;
else reg_24232921_result_delayed_u0<=reg_24232921_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2a60e877_u0<=1'h0;
else reg_2a60e877_u0<=reg_39c815b1_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1c7bd8c5_result_delayed_u0<=1'h0;
else reg_1c7bd8c5_result_delayed_u0<=reg_1c7bd8c5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_05b030d6_result_delayed_u0<=1'h0;
else reg_05b030d6_result_delayed_u0<=reg_05b030d6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6df7e814_result_delayed_u0<=1'h0;
else reg_6df7e814_result_delayed_u0<=reg_6df7e814_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0530331a_u0<=1'h0;
else reg_0530331a_u0<=reg_04a57b8c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5df79fda_u0<=1'h0;
else reg_5df79fda_u0<=reg_77668746_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2add40ec_u0<=1'h0;
else reg_2add40ec_u0<=reg_367fcb5d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_195de36c_u0<=1'h0;
else reg_195de36c_u0<=reg_710f71fd_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4f367a8e_result_delayed_u0<=1'h0;
else reg_4f367a8e_result_delayed_u0<=reg_4f367a8e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_70b8aa8a_u0<=1'h0;
else reg_70b8aa8a_u0<=reg_0b769204_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_52bc0089_u0<=1'h0;
else reg_52bc0089_u0<=reg_6dec38b5_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0fa7db18_result_delayed_result_delayed_u0<=1'h0;
else reg_0fa7db18_result_delayed_result_delayed_u0<=reg_0fa7db18_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_62bcd2be_result_delayed_result_delayed_u0<=1'h0;
else reg_62bcd2be_result_delayed_result_delayed_u0<=reg_62bcd2be_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01a00b9a_u0<=1'h0;
else reg_01a00b9a_u0<=reg_441fe928_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_08eb52d0_u0<=1'h0;
else reg_08eb52d0_u0<=reg_0f726638_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_68801c52_result_delayed_result_delayed_u0<=1'h0;
else reg_68801c52_result_delayed_result_delayed_u0<=reg_68801c52_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_66565274_result_delayed_u0<=1'h0;
else reg_66565274_result_delayed_u0<=reg_66565274_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3c2e9ca2_result_delayed_u0<=1'h0;
else reg_3c2e9ca2_result_delayed_u0<=reg_3c2e9ca2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5874fe30_u0<=1'h0;
else reg_5874fe30_u0<=reg_7bd0a7f4_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3a9ed8da_u0<=1'h0;
else reg_3a9ed8da_u0<=reg_4df0fb45_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6f2cfbe7_result_delayed_result_delayed_u0<=1'h0;
else reg_6f2cfbe7_result_delayed_result_delayed_u0<=reg_6f2cfbe7_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_24a21cbf_result_delayed_result_delayed_u0<=1'h0;
else reg_24a21cbf_result_delayed_result_delayed_u0<=reg_24a21cbf_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7ffc667d_result_delayed_result_delayed_u0<=1'h0;
else reg_7ffc667d_result_delayed_result_delayed_u0<=reg_7ffc667d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2efcd75c_result_delayed_u0<=1'h0;
else reg_2efcd75c_result_delayed_u0<=reg_2efcd75c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1796d9d9_u0<=1'h0;
else reg_1796d9d9_u0<=reg_52bc0089_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_58a2a0e3_result_delayed_u0<=1'h0;
else reg_58a2a0e3_result_delayed_u0<=reg_58a2a0e3_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_04da25b8_result_delayed_u0<=1'h0;
else reg_04da25b8_result_delayed_u0<=reg_04da25b8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00246672_u0<=1'h0;
else reg_00246672_u0<=reg_05b030d6_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6ec6926a_result_delayed_u0<=1'h0;
else reg_6ec6926a_result_delayed_u0<=reg_6ec6926a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_32c8d37c_result_delayed_u0<=1'h0;
else reg_32c8d37c_result_delayed_u0<=reg_32c8d37c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0b8053fe_result_delayed_result_delayed_u0<=1'h0;
else reg_0b8053fe_result_delayed_result_delayed_u0<=reg_0b8053fe_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0ee3ba53_result_delayed_result_delayed_u0<=1'h0;
else reg_0ee3ba53_result_delayed_result_delayed_u0<=reg_0ee3ba53_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2976ab2a_u0<=1'h0;
else reg_2976ab2a_u0<=reg_1098e4cf_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1fa5ca42_result_delayed_u0<=1'h0;
else reg_1fa5ca42_result_delayed_u0<=reg_1fa5ca42_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1457ec7b_result_delayed_u0<=1'h0;
else reg_1457ec7b_result_delayed_u0<=reg_1457ec7b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_68d00eb5_u0<=1'h0;
else reg_68d00eb5_u0<=reg_710efd1b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_68ca4866_result_delayed_u0<=1'h0;
else reg_68ca4866_result_delayed_u0<=reg_68ca4866_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_39c815b1_result_delayed_u0<=1'h0;
else reg_39c815b1_result_delayed_u0<=reg_39c815b1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1623704a_u0<=1'h0;
else reg_1623704a_u0<=reg_68e2082a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5451da38_u0<=1'h0;
else reg_5451da38_u0<=reg_640f5a91_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7d510c70_result_delayed_u0<=1'h0;
else reg_7d510c70_result_delayed_u0<=reg_7d510c70_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1036257e_result_delayed_u0<=1'h0;
else reg_1036257e_result_delayed_u0<=reg_1036257e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_18e93e99_u0<=1'h0;
else reg_18e93e99_u0<=reg_201eb03b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7999bbe8_u0<=1'h0;
else reg_7999bbe8_u0<=reg_4c7e6a09_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1418995e_result_delayed_u0<=1'h0;
else reg_1418995e_result_delayed_u0<=reg_1418995e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_677157b7_result_delayed_u0<=1'h0;
else reg_677157b7_result_delayed_u0<=reg_677157b7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4c7e6a09_u0<=1'h0;
else reg_4c7e6a09_u0<=reg_6f9e56f4_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_53090f63_result_delayed_u0<=1'h0;
else reg_53090f63_result_delayed_u0<=reg_53090f63_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_05b030d6_result_delayed_result_delayed_u0<=1'h0;
else reg_05b030d6_result_delayed_result_delayed_u0<=reg_05b030d6_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4235f44a_u0<=1'h0;
else reg_4235f44a_u0<=reg_26133792_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_142b80f2_result_delayed_u0<=1'h0;
else reg_142b80f2_result_delayed_u0<=reg_142b80f2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_09e28b61_u0<=1'h0;
else reg_09e28b61_u0<=reg_68801c52_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_227958fa_u0<=1'h0;
else reg_227958fa_u0<=reg_1fa5ca42_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_06efce9a_result_delayed_result_delayed_u0<=1'h0;
else reg_06efce9a_result_delayed_result_delayed_u0<=reg_06efce9a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_52bc0089_result_delayed_u0<=1'h0;
else reg_52bc0089_result_delayed_u0<=reg_52bc0089_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4e1c133b_result_delayed_result_delayed_u0<=1'h0;
else reg_4e1c133b_result_delayed_result_delayed_u0<=reg_4e1c133b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6028598b_result_delayed_result_delayed_u0<=1'h0;
else reg_6028598b_result_delayed_result_delayed_u0<=reg_6028598b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7bd0a7f4_result_delayed_u0<=1'h0;
else reg_7bd0a7f4_result_delayed_u0<=reg_7bd0a7f4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4d3893b7_u0<=1'h0;
else reg_4d3893b7_u0<=reg_747c90de_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4235f44a_result_delayed_u0<=1'h0;
else reg_4235f44a_result_delayed_u0<=reg_4235f44a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_690deb9c_u0<=1'h0;
else reg_690deb9c_u0<=reg_229d1ee4_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1ea77ba6_result_delayed_u0<=1'h0;
else reg_1ea77ba6_result_delayed_u0<=reg_1ea77ba6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1418995e_result_delayed_result_delayed_u0<=1'h0;
else reg_1418995e_result_delayed_result_delayed_u0<=reg_1418995e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_18ff3a6a_u0<=1'h0;
else reg_18ff3a6a_u0<=reg_1dd4f561_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2ed4804d_u0<=1'h0;
else reg_2ed4804d_u0<=reg_5674bffb_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_39c815b1_result_delayed_result_delayed_u0<=1'h0;
else reg_39c815b1_result_delayed_result_delayed_u0<=reg_39c815b1_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_640f5a91_u0<=1'h0;
else reg_640f5a91_u0<=reg_00af20e1_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1ad50076_u0<=1'h0;
else reg_1ad50076_u0<=reg_68ca4866_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1c1149c7_result_delayed_u0<=1'h0;
else reg_1c1149c7_result_delayed_u0<=reg_1c1149c7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4cc74cbd_result_delayed_result_delayed_u0<=1'h0;
else reg_4cc74cbd_result_delayed_result_delayed_u0<=reg_4cc74cbd_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0f726638_result_delayed_u0<=1'h0;
else reg_0f726638_result_delayed_u0<=reg_0f726638_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0a3ee092_u0<=1'h0;
else reg_0a3ee092_u0<=reg_4769eae6_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5451da38_result_delayed_u0<=1'h0;
else reg_5451da38_result_delayed_u0<=reg_5451da38_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1fa5ca42_result_delayed_result_delayed_u0<=1'h0;
else reg_1fa5ca42_result_delayed_result_delayed_u0<=reg_1fa5ca42_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4df0fb45_u0<=1'h0;
else reg_4df0fb45_u0<=reg_445ccdaa_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6092b844_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_6092b844_result_delayed_result_delayed_result_delayed_u0<=reg_6092b844_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_64049807_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_64049807_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_64049807_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_258244c0_result_delayed_u0<=1'h0;
else reg_258244c0_result_delayed_u0<=reg_258244c0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1457ec7b_result_delayed_result_delayed_u0<=1'h0;
else reg_1457ec7b_result_delayed_result_delayed_u0<=reg_1457ec7b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0b8053fe_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_0b8053fe_result_delayed_result_delayed_result_delayed_u0<=reg_0b8053fe_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1a0fb632_result_delayed_result_delayed_u0<=1'h0;
else reg_1a0fb632_result_delayed_result_delayed_u0<=reg_1a0fb632_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3c2e9ca2_result_delayed_result_delayed_u0<=1'h0;
else reg_3c2e9ca2_result_delayed_result_delayed_u0<=reg_3c2e9ca2_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0076a506_result_delayed_u0<=1'h0;
else reg_0076a506_result_delayed_u0<=reg_0076a506_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_75fb999e_result_delayed_u0<=1'h0;
else reg_75fb999e_result_delayed_u0<=reg_75fb999e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_15c73839_result_delayed_u0<=1'h0;
else reg_15c73839_result_delayed_u0<=reg_15c73839_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2f2401f0_u0<=1'h0;
else reg_2f2401f0_u0<=reg_7999bbe8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4235f44a_result_delayed_result_delayed_u0<=1'h0;
else reg_4235f44a_result_delayed_result_delayed_u0<=reg_4235f44a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_576a3720_result_delayed_u0<=1'h0;
else reg_576a3720_result_delayed_u0<=reg_576a3720_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7723f5fb_u0<=1'h0;
else reg_7723f5fb_u0<=reg_7807eb12_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_426d8380_result_delayed_u0<=1'h0;
else reg_426d8380_result_delayed_u0<=reg_426d8380_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_26133792_result_delayed_u0<=1'h0;
else reg_26133792_result_delayed_u0<=reg_26133792_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4d3893b7_result_delayed_u0<=1'h0;
else reg_4d3893b7_result_delayed_u0<=reg_4d3893b7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_228ef2dc_result_delayed_u0<=1'h0;
else reg_228ef2dc_result_delayed_u0<=reg_228ef2dc_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_43da3530_u0<=1'h0;
else reg_43da3530_u0<=reg_4235f44a_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_22603c8b_u0<=1'h0;
else reg_22603c8b_u0<=reg_343e0093_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_21c538b9_result_delayed_u0<=1'h0;
else reg_21c538b9_result_delayed_u0<=reg_21c538b9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_677157b7_result_delayed_result_delayed_u0<=1'h0;
else reg_677157b7_result_delayed_result_delayed_u0<=reg_677157b7_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_576a3720_result_delayed_result_delayed_u0<=1'h0;
else reg_576a3720_result_delayed_result_delayed_u0<=reg_576a3720_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_304f02b2_u0<=1'h0;
else reg_304f02b2_u0<=reg_426d8380_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0986382d_result_delayed_u0<=1'h0;
else reg_0986382d_result_delayed_u0<=reg_0986382d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6d17e172_result_delayed_u0<=1'h0;
else reg_6d17e172_result_delayed_u0<=reg_6d17e172_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_735b3058_u0<=1'h0;
else reg_735b3058_u0<=reg_36ce22d8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_24a21cbf_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_24a21cbf_result_delayed_result_delayed_result_delayed_u0<=reg_24a21cbf_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_201eb03b_result_delayed_u0<=1'h0;
else reg_201eb03b_result_delayed_u0<=reg_201eb03b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0bcf08c6_u0<=1'h0;
else reg_0bcf08c6_u0<=reg_070292d1_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_747c90de_result_delayed_result_delayed_u0<=1'h0;
else reg_747c90de_result_delayed_result_delayed_u0<=reg_747c90de_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0a6a1b0e_result_delayed_u0<=1'h0;
else reg_0a6a1b0e_result_delayed_u0<=reg_0a6a1b0e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2f9dd090_u0<=1'h0;
else reg_2f9dd090_u0<=reg_7d231906_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_30e8bfe6_u0<=1'h0;
else reg_30e8bfe6_u0<=reg_180dc380_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_445ccdaa_result_delayed_u0<=1'h0;
else reg_445ccdaa_result_delayed_u0<=reg_445ccdaa_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_55edd085_result_delayed_u0<=1'h0;
else reg_55edd085_result_delayed_u0<=reg_55edd085_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7807eb12_u0<=1'h0;
else reg_7807eb12_u0<=reg_4ffb5ab4_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1098e4cf_result_delayed_u0<=1'h0;
else reg_1098e4cf_result_delayed_u0<=reg_1098e4cf_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_242facb3_result_delayed_result_delayed_u0<=1'h0;
else reg_242facb3_result_delayed_result_delayed_u0<=reg_242facb3_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_77d7ef15_result_delayed_result_delayed_u0<=1'h0;
else reg_77d7ef15_result_delayed_result_delayed_u0<=reg_77d7ef15_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7723f5fb_result_delayed_u0<=1'h0;
else reg_7723f5fb_result_delayed_u0<=reg_7723f5fb_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0b769204_result_delayed_u0<=1'h0;
else reg_0b769204_result_delayed_u0<=reg_0b769204_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_367fcb5d_result_delayed_u0<=1'h0;
else reg_367fcb5d_result_delayed_u0<=reg_367fcb5d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_387904fe_result_delayed_u0<=1'h0;
else reg_387904fe_result_delayed_u0<=reg_387904fe_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_104b8d92_result_delayed_u0<=1'h0;
else reg_104b8d92_result_delayed_u0<=reg_104b8d92_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2537f8df_result_delayed_u0<=1'h0;
else reg_2537f8df_result_delayed_u0<=reg_2537f8df_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_04a57b8c_u0<=1'h0;
else reg_04a57b8c_u0<=reg_64daf8c4_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2f9dd090_result_delayed_u0<=1'h0;
else reg_2f9dd090_result_delayed_u0<=reg_2f9dd090_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7d61464a_u0<=1'h0;
else reg_7d61464a_u0<=reg_6a79fa17_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4235f44a_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_4235f44a_result_delayed_result_delayed_result_delayed_u0<=reg_4235f44a_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_343e0093_result_delayed_u0<=1'h0;
else reg_343e0093_result_delayed_u0<=reg_343e0093_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_77668746_result_delayed_result_delayed_u0<=1'h0;
else reg_77668746_result_delayed_result_delayed_u0<=reg_77668746_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00af20e1_result_delayed_u0<=1'h0;
else reg_00af20e1_result_delayed_u0<=reg_00af20e1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_35c4a85b_result_delayed_u0<=1'h0;
else reg_35c4a85b_result_delayed_u0<=reg_35c4a85b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_64daf8c4_result_delayed_u0<=1'h0;
else reg_64daf8c4_result_delayed_u0<=reg_64daf8c4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_18ad0cb7_result_delayed_u0<=1'h0;
else reg_18ad0cb7_result_delayed_u0<=reg_18ad0cb7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_68801c52_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_68801c52_result_delayed_result_delayed_result_delayed_u0<=reg_68801c52_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_49242595_result_delayed_u0<=1'h0;
else reg_49242595_result_delayed_u0<=reg_49242595_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1680ee34_result_delayed_u0<=1'h0;
else reg_1680ee34_result_delayed_u0<=reg_1680ee34_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2c8dcfcc_u0<=1'h0;
else reg_2c8dcfcc_u0<=reg_5650d91a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_54ef10cf_result_delayed_u0<=1'h0;
else reg_54ef10cf_result_delayed_u0<=reg_54ef10cf_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_35d48481_result_delayed_u0<=1'h0;
else reg_35d48481_result_delayed_u0<=reg_35d48481_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_36ce22d8_result_delayed_u0<=1'h0;
else reg_36ce22d8_result_delayed_u0<=reg_36ce22d8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0425c0a1_result_delayed_u0<=1'h0;
else reg_0425c0a1_result_delayed_u0<=reg_0425c0a1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4a77e6f2_result_delayed_u0<=1'h0;
else reg_4a77e6f2_result_delayed_u0<=reg_4a77e6f2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5650d91a_u0<=1'h0;
else reg_5650d91a_u0<=reg_32c8d37c_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_796241e6_result_delayed_u0<=1'h0;
else reg_796241e6_result_delayed_u0<=reg_796241e6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_08eb52d0_result_delayed_u0<=1'h0;
else reg_08eb52d0_result_delayed_u0<=reg_08eb52d0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6a79fa17_result_delayed_u0<=1'h0;
else reg_6a79fa17_result_delayed_u0<=reg_6a79fa17_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_32a37dec_u0<=1'h0;
else reg_32a37dec_u0<=reg_2a321227_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_38d95389_u0<=1'h0;
else reg_38d95389_u0<=reg_6bf613ee_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_70b8aa8a_result_delayed_u0<=1'h0;
else reg_70b8aa8a_result_delayed_u0<=reg_70b8aa8a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_44a5d7f1_u0<=1'h0;
else reg_44a5d7f1_u0<=reg_00246672_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5674bffb_result_delayed_u0<=1'h0;
else reg_5674bffb_result_delayed_u0<=reg_5674bffb_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4769eae6_result_delayed_u0<=1'h0;
else reg_4769eae6_result_delayed_u0<=reg_4769eae6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4ffb5ab4_result_delayed_result_delayed_u0<=1'h0;
else reg_4ffb5ab4_result_delayed_result_delayed_u0<=reg_4ffb5ab4_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_441fe928_result_delayed_u0<=1'h0;
else reg_441fe928_result_delayed_u0<=reg_441fe928_u0;
end
assign and_u2220_u0=and_u2214_u0&and_u2222_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0a6a1b0e_result_delayed_result_delayed_u0<=1'h0;
else reg_0a6a1b0e_result_delayed_result_delayed_u0<=reg_0a6a1b0e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6bf613ee_result_delayed_u0<=1'h0;
else reg_6bf613ee_result_delayed_u0<=reg_6bf613ee_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_710efd1b_result_delayed_u0<=1'h0;
else reg_710efd1b_result_delayed_u0<=reg_710efd1b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1dd4f561_result_delayed_result_delayed_u0<=1'h0;
else reg_1dd4f561_result_delayed_result_delayed_u0<=reg_1dd4f561_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_09302a5b_u0<=1'h0;
else reg_09302a5b_u0<=reg_2c8dcfcc_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_18e93e99_result_delayed_u0<=1'h0;
else reg_18e93e99_result_delayed_u0<=reg_18e93e99_u0;
end
assign or_u690_u0=and_u2220_u0|and_u2218_u0;
assign mux_u224=(and_u2220_u0)?1'h1:1'h0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0b8053fe_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_0b8053fe_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_0b8053fe_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_70b8aa8a_result_delayed_result_delayed_u0<=1'h0;
else reg_70b8aa8a_result_delayed_result_delayed_u0<=reg_70b8aa8a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_227958fa_result_delayed_u0<=1'h0;
else reg_227958fa_result_delayed_u0<=reg_227958fa_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_382aec0c_result_delayed_result_delayed_u0<=1'h0;
else reg_382aec0c_result_delayed_result_delayed_u0<=reg_382aec0c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0fa7db18_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_0fa7db18_result_delayed_result_delayed_result_delayed_u0<=reg_0fa7db18_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_09408e3d_u0<=1'h0;
else reg_09408e3d_u0<=reg_39d6e99f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6092b844_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_6092b844_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_6092b844_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4bbdc680_result_delayed_u0<=1'h0;
else reg_4bbdc680_result_delayed_u0<=reg_4bbdc680_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_13cde2f7_result_delayed_u0<=1'h0;
else reg_13cde2f7_result_delayed_u0<=reg_13cde2f7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_343e0093_result_delayed_result_delayed_u0<=1'h0;
else reg_343e0093_result_delayed_result_delayed_u0<=reg_343e0093_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7999bbe8_result_delayed_u0<=1'h0;
else reg_7999bbe8_result_delayed_u0<=reg_7999bbe8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4e289baa_result_delayed_u0<=1'h0;
else reg_4e289baa_result_delayed_u0<=reg_4e289baa_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1a79d7d6_result_delayed_u0<=1'h0;
else reg_1a79d7d6_result_delayed_u0<=reg_1a79d7d6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1dd4f561_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_1dd4f561_result_delayed_result_delayed_result_delayed_u0<=reg_1dd4f561_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1a837eb0_result_delayed_u0<=1'h0;
else reg_1a837eb0_result_delayed_u0<=reg_1a837eb0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7bfae876_u0<=1'h0;
else reg_7bfae876_u0<=reg_5bc0cf31_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7d46a529_result_delayed_u0<=1'h0;
else reg_7d46a529_result_delayed_u0<=reg_7d46a529_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_180dc380_u0<=1'h0;
else reg_180dc380_u0<=reg_6df7e814_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3a9ed8da_result_delayed_u0<=1'h0;
else reg_3a9ed8da_result_delayed_u0<=reg_3a9ed8da_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_70b8aa8a_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_70b8aa8a_result_delayed_result_delayed_result_delayed_u0<=reg_70b8aa8a_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_32c8d37c_result_delayed_result_delayed_u0<=1'h0;
else reg_32c8d37c_result_delayed_result_delayed_u0<=reg_32c8d37c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_64789d0a_result_delayed_u0<=1'h0;
else reg_64789d0a_result_delayed_u0<=reg_64789d0a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_42536b9e_result_delayed_u0<=1'h0;
else reg_42536b9e_result_delayed_u0<=reg_42536b9e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_229d1ee4_result_delayed_result_delayed_u0<=1'h0;
else reg_229d1ee4_result_delayed_result_delayed_u0<=reg_229d1ee4_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1cd8b4df_result_delayed_u0<=1'h0;
else reg_1cd8b4df_result_delayed_u0<=reg_1cd8b4df_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_06dc9aa2_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_06dc9aa2_result_delayed_result_delayed_result_delayed_u0<=reg_06dc9aa2_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6f9e56f4_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_6f9e56f4_result_delayed_result_delayed_result_delayed_u0<=reg_6f9e56f4_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_304f02b2_result_delayed_u0<=1'h0;
else reg_304f02b2_result_delayed_u0<=reg_304f02b2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5ee7823f_result_delayed_u0<=1'h0;
else reg_5ee7823f_result_delayed_u0<=reg_5ee7823f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6df7e814_result_delayed_result_delayed_u0<=1'h0;
else reg_6df7e814_result_delayed_result_delayed_u0<=reg_6df7e814_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4a5adf10_result_delayed_result_delayed_u0<=1'h0;
else reg_4a5adf10_result_delayed_result_delayed_u0<=reg_4a5adf10_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_18ff3a6a_result_delayed_u0<=1'h0;
else reg_18ff3a6a_result_delayed_u0<=reg_18ff3a6a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4ffb5ab4_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_4ffb5ab4_result_delayed_result_delayed_result_delayed_u0<=reg_4ffb5ab4_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5e4d335d_result_delayed_result_delayed_u0<=1'h0;
else reg_5e4d335d_result_delayed_result_delayed_u0<=reg_5e4d335d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_528f4535_u0<=1'h0;
else reg_528f4535_u0<=reg_76ad5fc6_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_242facb3_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_242facb3_result_delayed_result_delayed_result_delayed_u0<=reg_242facb3_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00246672_result_delayed_u0<=1'h0;
else reg_00246672_result_delayed_u0<=reg_00246672_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_10810426_result_delayed_u0<=1'h0;
else reg_10810426_result_delayed_u0<=reg_10810426_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_09e28b61_result_delayed_u0<=1'h0;
else reg_09e28b61_result_delayed_u0<=reg_09e28b61_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a05baae_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_7a05baae_result_delayed_result_delayed_result_delayed_u0<=reg_7a05baae_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0f5456f1_result_delayed_u0<=1'h0;
else reg_0f5456f1_result_delayed_u0<=reg_0f5456f1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_710f71fd_result_delayed_result_delayed_u0<=1'h0;
else reg_710f71fd_result_delayed_result_delayed_u0<=reg_710f71fd_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_426d8380_result_delayed_result_delayed_u0<=1'h0;
else reg_426d8380_result_delayed_result_delayed_u0<=reg_426d8380_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6d759d56_result_delayed_result_delayed_u0<=1'h0;
else reg_6d759d56_result_delayed_result_delayed_u0<=reg_6d759d56_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_09e28b61_result_delayed_result_delayed_u0<=1'h0;
else reg_09e28b61_result_delayed_result_delayed_u0<=reg_09e28b61_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_640dac03_result_delayed_u0<=1'h0;
else reg_640dac03_result_delayed_u0<=reg_640dac03_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2a321227_result_delayed_u0<=1'h0;
else reg_2a321227_result_delayed_u0<=reg_2a321227_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2c8dcfcc_result_delayed_u0<=1'h0;
else reg_2c8dcfcc_result_delayed_u0<=reg_2c8dcfcc_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6dec38b5_result_delayed_u0<=1'h0;
else reg_6dec38b5_result_delayed_u0<=reg_6dec38b5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5bc0cf31_result_delayed_result_delayed_u0<=1'h0;
else reg_5bc0cf31_result_delayed_result_delayed_u0<=reg_5bc0cf31_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_02369e1a_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_02369e1a_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_02369e1a_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_424e119f_u0<=1'h0;
else reg_424e119f_u0<=reg_405c3132_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5c7b4c7d_result_delayed_result_delayed_u0<=1'h0;
else reg_5c7b4c7d_result_delayed_result_delayed_u0<=reg_5c7b4c7d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_070292d1_result_delayed_u0<=1'h0;
else reg_070292d1_result_delayed_u0<=reg_070292d1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7e3e122c_result_delayed_u0<=1'h0;
else reg_7e3e122c_result_delayed_u0<=reg_7e3e122c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_05b030d6_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_05b030d6_result_delayed_result_delayed_result_delayed_u0<=reg_05b030d6_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_405c3132_result_delayed_u0<=1'h0;
else reg_405c3132_result_delayed_u0<=reg_405c3132_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4a77e6f2_result_delayed_result_delayed_u0<=1'h0;
else reg_4a77e6f2_result_delayed_result_delayed_u0<=reg_4a77e6f2_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0b38372d_result_delayed_result_delayed_u0<=1'h0;
else reg_0b38372d_result_delayed_result_delayed_u0<=reg_0b38372d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0d9b29cf_result_delayed_u0<=1'h0;
else reg_0d9b29cf_result_delayed_u0<=reg_0d9b29cf_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5ee7823f_result_delayed_result_delayed_u0<=1'h0;
else reg_5ee7823f_result_delayed_result_delayed_u0<=reg_5ee7823f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2f9dd090_result_delayed_result_delayed_u0<=1'h0;
else reg_2f9dd090_result_delayed_result_delayed_u0<=reg_2f9dd090_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1098e4cf_result_delayed_result_delayed_u0<=1'h0;
else reg_1098e4cf_result_delayed_result_delayed_u0<=reg_1098e4cf_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_39d6e99f_result_delayed_u0<=1'h0;
else reg_39d6e99f_result_delayed_u0<=reg_39d6e99f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7d231906_result_delayed_u0<=1'h0;
else reg_7d231906_result_delayed_u0<=reg_7d231906_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_47aed7f7_result_delayed_u0<=1'h0;
else reg_47aed7f7_result_delayed_u0<=reg_47aed7f7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_104b8d92_result_delayed_result_delayed_u0<=1'h0;
else reg_104b8d92_result_delayed_result_delayed_u0<=reg_104b8d92_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1dce6126_result_delayed_u0<=1'h0;
else reg_1dce6126_result_delayed_u0<=reg_1dce6126_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_183f91d8_result_delayed_u0<=1'h0;
else reg_183f91d8_result_delayed_u0<=reg_183f91d8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_68e2082a_result_delayed_u0<=1'h0;
else reg_68e2082a_result_delayed_u0<=reg_68e2082a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_64daf8c4_result_delayed_result_delayed_u0<=1'h0;
else reg_64daf8c4_result_delayed_result_delayed_u0<=reg_64daf8c4_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_76ad5fc6_result_delayed_u0<=1'h0;
else reg_76ad5fc6_result_delayed_u0<=reg_76ad5fc6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_06efce9a_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_06efce9a_result_delayed_result_delayed_result_delayed_u0<=reg_06efce9a_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6dec38b5_result_delayed_result_delayed_u0<=1'h0;
else reg_6dec38b5_result_delayed_result_delayed_u0<=reg_6dec38b5_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_68ca4866_result_delayed_result_delayed_u0<=1'h0;
else reg_68ca4866_result_delayed_result_delayed_u0<=reg_68ca4866_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2efcd75c_result_delayed_result_delayed_u0<=1'h0;
else reg_2efcd75c_result_delayed_result_delayed_u0<=reg_2efcd75c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6320b243_result_delayed_result_delayed_u0<=1'h0;
else reg_6320b243_result_delayed_result_delayed_u0<=reg_6320b243_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2d8f78b3_result_delayed_u0<=1'h0;
else reg_2d8f78b3_result_delayed_u0<=reg_2d8f78b3_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0f7cf45c_u0<=1'h0;
else reg_0f7cf45c_u0<=and_u2221_u0;
end
assign or_u691_u0=and_u2221_u0|and_u2220_u0;
assign mux_u225_u0=(and_u2221_u0)?32'h4:32'h200;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0f7cf45c_result_delayed_u0<=1'h0;
else reg_0f7cf45c_result_delayed_u0<=reg_0f7cf45c_u0;
end
assign or_u692_u0=and_u2221_u0|and_u2220_u0;
assign or_u693_u0=and_u2221_u0|and_u2220_u0;
assign and_u2221_u0=and_u2213_u0&and_u2223_u0;
assign or_u694_u0=reg_1f5cf7c4_result_delayed_u0|or_u689_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1f5cf7c4_u0<=1'h0;
else reg_1f5cf7c4_u0<=reg_0f7cf45c_result_delayed_result_delayed_u0;
end
assign and_u2222_u0=and_u2212_u0&and_u2223_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1f5cf7c4_result_delayed_u0<=1'h0;
else reg_1f5cf7c4_result_delayed_u0<=reg_1f5cf7c4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0f7cf45c_result_delayed_result_delayed_u0<=1'h0;
else reg_0f7cf45c_result_delayed_result_delayed_u0<=reg_0f7cf45c_result_delayed_u0;
end
assign or_u695_u0=and_u2221_u0|and_u2220_u0;
assign mux_u226_u0=(and_u2221_u0)?1'h1:mux_u224;
assign or_u696_u0=and_u2221_u0|or_u690_u0;
assign and_u2223_u0=and_u2211_u0&and_u2242_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1769529a_u0<=1'h0;
else reg_1769529a_u0<=and_u2224_u0;
end
assign or_u697_u0=or_u694_u0|reg_1769529a_u0;
assign and_u2224_u0=and_u2210_u0&and_u2242_u0;
assign equals_u118_a_signed={31'b0, port_768be70f_};
assign equals_u118_b_signed=32'h1;
assign equals_u118=equals_u118_a_signed==equals_u118_b_signed;
assign and_u2225_u0=and_u2242_u0&equals_u118;
assign and_u2226_u0=and_u2242_u0&not_u409_u0;
assign not_u409_u0=~equals_u118;
assign not_u410_u0=~port_607140ed_;
assign and_u2227_u0=and_u2241_u0&port_607140ed_;
assign and_u2228_u0=and_u2241_u0&not_u410_u0;
assign lessThan_u51_a_signed=port_30496c3f_;
assign lessThan_u51_b_signed=port_1bf015b7_;
assign lessThan_u51=lessThan_u51_a_signed<lessThan_u51_b_signed;
assign not_u411_u0=~lessThan_u51;
assign and_u2229_u0=and_u2238_u0&not_u411_u0;
assign and_u2230_u0=and_u2238_u0&lessThan_u51;
assign and_u2231_u0=and_u2236_u0&port_6a29d19a_;
assign not_u412_u0=~port_6a29d19a_;
assign and_u2232_u0=and_u2236_u0&not_u412_u0;
assign add=port_30496c3f_+32'h0;
assign and_u2233_u0=and_u2235_u0&port_4a47b2ff_;
assign simplePinWrite_u368=and_u2235_u0&{1{and_u2235_u0}};
assign simplePinWrite_u369=port_7dc406cd_;
assign simplePinWrite_u370=16'h1&{16{1'h1}};
assign add_u167=port_30496c3f_+32'h1;
always @(posedge CLK)
begin
if (and_u2235_u0)
syncEnable_u317<=port_7dc406cd_;
end
assign mux_u227_u0=(reg_3543084e_u0)?syncEnable_u317:syncEnable_u318_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3543084e_u0<=1'h0;
else reg_3543084e_u0<=and_u2235_u0;
end
assign and_u2234_u0=and_u2232_u0&and_u2236_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u145<=1'h0;
else and_delayed_u145<=and_u2234_u0;
end
always @(posedge CLK)
begin
if (and_u2236_u0)
syncEnable_u318_u0<=mux_u238_u0;
end
assign and_u2235_u0=and_u2231_u0&and_u2236_u0;
always @(posedge CLK)
begin
if (and_u2238_u0)
syncEnable_u319_u0<=mux_u239_u0;
end
always @(posedge CLK)
begin
if (and_u2238_u0)
syncEnable_u320_u0<=mux_u238_u0;
end
assign mux_u228_u0=(reg_5a8744bc_u0)?syncEnable_u320_u0:mux_u227_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_394c9807_u0<=1'h0;
else reg_394c9807_u0<=and_u2236_u0;
end
assign mux_u229_u0=(reg_5a8744bc_u0)?32'h0:syncEnable_u319_u0;
assign and_u2236_u0=and_u2230_u0&and_u2238_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5a8744bc_u0<=1'h0;
else reg_5a8744bc_u0<=and_u2237_u0;
end
assign and_u2237_u0=and_u2229_u0&and_u2238_u0;
assign mux_u230_u0=(reg_371d79bc_u0)?syncEnable_u321_u0:mux_u229_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_371d79bc_u0<=1'h0;
else reg_371d79bc_u0<=and_u2239_u0;
end
assign and_u2238_u0=and_u2227_u0&and_u2241_u0;
always @(posedge CLK)
begin
if (and_u2241_u0)
syncEnable_u321_u0<=mux_u239_u0;
end
assign and_u2239_u0=and_u2228_u0&and_u2241_u0;
always @(posedge CLK)
begin
if (and_u2241_u0)
syncEnable_u322_u0<=mux_u238_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u146_u0<=1'h0;
else and_delayed_u146_u0<=and_u2238_u0;
end
assign mux_u231_u0=(reg_371d79bc_u0)?syncEnable_u322_u0:mux_u228_u0;
assign mux_u232_u0=(and_delayed_u148_u0)?mux_u230_u0:syncEnable_u324_u0;
assign and_u2240_u0=and_u2226_u0&and_u2242_u0;
assign and_u2241_u0=and_u2225_u0&and_u2242_u0;
assign mux_u233_u0=(and_delayed_u148_u0)?mux_u231_u0:syncEnable_u323_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u147_u0<=1'h0;
else and_delayed_u147_u0<=and_u2240_u0;
end
always @(posedge CLK)
begin
if (and_u2242_u0)
syncEnable_u323_u0<=mux_u238_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u148_u0<=1'h0;
else and_delayed_u148_u0<=and_u2241_u0;
end
always @(posedge CLK)
begin
if (and_u2242_u0)
syncEnable_u324_u0<=mux_u239_u0;
end
assign mux_u234_u0=(or_u695_u0)?32'h0:add_u167;
assign or_u698_u0=or_u695_u0|and_u2235_u0;
assign or_u699_u0=or_u692_u0|and_u2237_u0;
assign mux_u235_u0=(or_u692_u0)?1'h1:1'h0;
assign mux_u236_u0=(or_u696_u0)?mux_u226_u0:1'h0;
assign or_u700_u0=or_u696_u0|and_u2237_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
block_GO_delayed_u8<=1'h0;
else block_GO_delayed_u8<=and_u2242_u0;
end
always @(posedge CLK)
begin
if (block_GO_delayed_u8)
latch_2c039393_reg<=mux_u233_u0;
end
assign latch_2c039393_out=(block_GO_delayed_u8)?mux_u233_u0:latch_2c039393_reg;
always @(posedge CLK)
begin
if (block_GO_delayed_u8)
latch_36791ce1_reg<=mux_u232_u0;
end
assign latch_36791ce1_out=(block_GO_delayed_u8)?mux_u232_u0:latch_36791ce1_reg;
assign mux_u237_u0=(or_u691_u0)?{22'b0, mux_u225_u0[9], 6'b0, mux_u225_u0[2], 2'b0}:32'hffffffff;
assign or_u701_u0=or_u691_u0|and_u2237_u0;
assign and_u2242_u0=or_u702_u0&or_u702_u0;
always @(posedge CLK)
begin
if (or_u697_u0)
fbReg_Out1Portvalue_u1<=latch_2c039393_out;
end
always @(posedge CLK)
begin
if (reg_01da6964_u0)
syncEnable_u325_u0<=RESET;
end
assign mux_u238_u0=(reg_01da6964_u0)?16'h0:fbReg_Out1Portvalue_u1;
assign or_u702_u0=reg_01da6964_u0|loopControl_u5;
always @(posedge CLK)
begin
if (or_u697_u0)
fbReg_temp_fsmOldState_resized_HH2_xy_4_u0<=latch_36791ce1_out;
end
assign mux_u239_u0=(reg_01da6964_u0)?32'h0:fbReg_temp_fsmOldState_resized_HH2_xy_4_u0;
always @(posedge CLK or posedge syncEnable_u325_u0)
begin
if (syncEnable_u325_u0)
loopControl_u5<=1'h0;
else loopControl_u5<=or_u697_u0;
end
assign or_u703_u0=GO|or_u693_u0;
assign or_u704_u0=GO|or_u700_u0;
assign mux_u240_u0=(GO)?1'h0:mux_u236_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01da6964_u0<=1'h0;
else reg_01da6964_u0<=reg_1c62611c_u0;
end
assign or_u705_u0=GO|or_u699_u0;
assign mux_u241_u0=(GO)?1'h0:mux_u235_u0;
assign or_u706_u0=GO|or_u701_u0;
assign mux_u242_u0=(GO)?32'hffffffff:mux_u237_u0;
assign or_u707_u0=GO|or_u698_u0;
assign mux_u243_u0=(GO)?32'h0:mux_u234_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1c62611c_u0<=1'h0;
else reg_1c62611c_u0<=GO;
end
assign RESULT=or_u703_u0;
assign RESULT_u1334=32'h0;
assign RESULT_u1335=or_u704_u0;
assign RESULT_u1336=mux_u240_u0;
assign RESULT_u1337=or_u707_u0;
assign RESULT_u1338=mux_u243_u0;
assign RESULT_u1339=or_u706_u0;
assign RESULT_u1340=mux_u242_u0;
assign RESULT_u1341=or_u705_u0;
assign RESULT_u1342=mux_u241_u0;
assign RESULT_u1343=and_u2235_u0;
assign RESULT_u1344=add;
assign RESULT_u1345=3'h1;
assign RESULT_u1346=simplePinWrite;
assign RESULT_u1347=simplePinWrite_u368;
assign RESULT_u1348=simplePinWrite_u366;
assign RESULT_u1349=simplePinWrite_u367;
assign RESULT_u1350=simplePinWrite_u370;
assign RESULT_u1351=simplePinWrite_u369;
assign DONE=1'h0;
endmodule



module resized_HH2_xy_endianswapper_20687a96_(endianswapper_20687a96_in, endianswapper_20687a96_out);
input	[31:0]	endianswapper_20687a96_in;
output	[31:0]	endianswapper_20687a96_out;
assign endianswapper_20687a96_out=endianswapper_20687a96_in;
endmodule



module resized_HH2_xy_endianswapper_56cc1fa2_(endianswapper_56cc1fa2_in, endianswapper_56cc1fa2_out);
input	[31:0]	endianswapper_56cc1fa2_in;
output	[31:0]	endianswapper_56cc1fa2_out;
assign endianswapper_56cc1fa2_out=endianswapper_56cc1fa2_in;
endmodule



module resized_HH2_xy_stateVar_Out1TokenIndex(bus_7ed6fa76_, bus_763548e3_, bus_51456afc_, bus_44270e5a_, bus_159d7a35_);
input		bus_7ed6fa76_;
input		bus_763548e3_;
input		bus_51456afc_;
input	[31:0]	bus_44270e5a_;
output	[31:0]	bus_159d7a35_;
reg	[31:0]	stateVar_Out1TokenIndex_u1=32'h0;
wire	[31:0]	endianswapper_20687a96_out;
wire	[31:0]	endianswapper_56cc1fa2_out;
always @(posedge bus_7ed6fa76_ or posedge bus_763548e3_)
begin
if (bus_763548e3_)
stateVar_Out1TokenIndex_u1<=32'h0;
else if (bus_51456afc_)
stateVar_Out1TokenIndex_u1<=endianswapper_20687a96_out;
end
assign bus_159d7a35_=endianswapper_56cc1fa2_out;
resized_HH2_xy_endianswapper_20687a96_ resized_HH2_xy_endianswapper_20687a96__1(.endianswapper_20687a96_in(bus_44270e5a_), 
  .endianswapper_20687a96_out(endianswapper_20687a96_out));
resized_HH2_xy_endianswapper_56cc1fa2_ resized_HH2_xy_endianswapper_56cc1fa2__1(.endianswapper_56cc1fa2_in(stateVar_Out1TokenIndex_u1), 
  .endianswapper_56cc1fa2_out(endianswapper_56cc1fa2_out));
endmodule



module resized_HH2_xy_forge_memory_512x16_23(CLK, EN, WE, ADDR, DIN, DOUT, DONE);
input		CLK;
input		EN;
input		WE;
input	[31:0]	ADDR;
input	[15:0]	DIN;
output	[15:0]	DOUT;
output		DONE;
wire		we_0;
wire	[15:0]	pre_dout_0;
wire		we_1;
wire	[15:0]	pre_dout_1;
wire		we_2;
wire	[15:0]	pre_dout_2;
wire		we_3;
wire	[15:0]	pre_dout_3;
reg	[15:0]	mux_out;
reg		wen_done;
assign we_0=WE&(ADDR[31:7]==25'h0);
assign we_1=WE&(ADDR[31:7]==25'h1);
assign we_2=WE&(ADDR[31:7]==25'h2);
assign we_3=WE&(ADDR[31:7]==25'h3);
always @(ADDR or pre_dout_0 or pre_dout_1 or pre_dout_2 or pre_dout_3)
begin
case (ADDR[31:7])25'd0:mux_out=pre_dout_0;
25'd1:mux_out=pre_dout_1;
25'd2:mux_out=pre_dout_2;
25'd3:mux_out=pre_dout_3;
default:mux_out=16'h0;
endcase end
always @(posedge CLK)
begin
wen_done<=WE;
end
assign DOUT=mux_out;
assign DONE=EN&!WE|wen_done;
//  Memory array element: COL: 0, ROW: 0
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_64(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[0]), .O(pre_dout_0[0]));
//  Memory array element: COL: 0, ROW: 1
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_65(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[1]), .O(pre_dout_0[1]));
//  Memory array element: COL: 0, ROW: 2
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_66(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[2]), .O(pre_dout_0[2]));
//  Memory array element: COL: 0, ROW: 3
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_67(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[3]), .O(pre_dout_0[3]));
//  Memory array element: COL: 0, ROW: 4
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_68(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[4]), .O(pre_dout_0[4]));
//  Memory array element: COL: 0, ROW: 5
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_69(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[5]), .O(pre_dout_0[5]));
//  Memory array element: COL: 0, ROW: 6
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_70(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[6]), .O(pre_dout_0[6]));
//  Memory array element: COL: 0, ROW: 7
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_71(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[7]), .O(pre_dout_0[7]));
//  Memory array element: COL: 0, ROW: 8
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_72(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[8]), .O(pre_dout_0[8]));
//  Memory array element: COL: 0, ROW: 9
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_73(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[9]), .O(pre_dout_0[9]));
//  Memory array element: COL: 0, ROW: 10
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_74(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[10]), .O(pre_dout_0[10]));
//  Memory array element: COL: 0, ROW: 11
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_75(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[11]), .O(pre_dout_0[11]));
//  Memory array element: COL: 0, ROW: 12
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_76(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[12]), .O(pre_dout_0[12]));
//  Memory array element: COL: 0, ROW: 13
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_77(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[13]), .O(pre_dout_0[13]));
//  Memory array element: COL: 0, ROW: 14
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_78(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[14]), .O(pre_dout_0[14]));
//  Memory array element: COL: 0, ROW: 15
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_79(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[15]), .O(pre_dout_0[15]));
//  Memory array element: COL: 1, ROW: 0
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_80(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[0]), .O(pre_dout_1[0]));
//  Memory array element: COL: 1, ROW: 1
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_81(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[1]), .O(pre_dout_1[1]));
//  Memory array element: COL: 1, ROW: 2
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_82(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[2]), .O(pre_dout_1[2]));
//  Memory array element: COL: 1, ROW: 3
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_83(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[3]), .O(pre_dout_1[3]));
//  Memory array element: COL: 1, ROW: 4
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_84(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[4]), .O(pre_dout_1[4]));
//  Memory array element: COL: 1, ROW: 5
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_85(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[5]), .O(pre_dout_1[5]));
//  Memory array element: COL: 1, ROW: 6
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_86(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[6]), .O(pre_dout_1[6]));
//  Memory array element: COL: 1, ROW: 7
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_87(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[7]), .O(pre_dout_1[7]));
//  Memory array element: COL: 1, ROW: 8
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_88(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[8]), .O(pre_dout_1[8]));
//  Memory array element: COL: 1, ROW: 9
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_89(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[9]), .O(pre_dout_1[9]));
//  Memory array element: COL: 1, ROW: 10
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_90(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[10]), .O(pre_dout_1[10]));
//  Memory array element: COL: 1, ROW: 11
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_91(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[11]), .O(pre_dout_1[11]));
//  Memory array element: COL: 1, ROW: 12
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_92(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[12]), .O(pre_dout_1[12]));
//  Memory array element: COL: 1, ROW: 13
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_93(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[13]), .O(pre_dout_1[13]));
//  Memory array element: COL: 1, ROW: 14
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_94(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[14]), .O(pre_dout_1[14]));
//  Memory array element: COL: 1, ROW: 15
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_95(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[15]), .O(pre_dout_1[15]));
//  Memory array element: COL: 2, ROW: 0
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_96(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[0]), .O(pre_dout_2[0]));
//  Memory array element: COL: 2, ROW: 1
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_97(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[1]), .O(pre_dout_2[1]));
//  Memory array element: COL: 2, ROW: 2
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_98(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[2]), .O(pre_dout_2[2]));
//  Memory array element: COL: 2, ROW: 3
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_99(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[3]), .O(pre_dout_2[3]));
//  Memory array element: COL: 2, ROW: 4
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_100(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[4]), .O(pre_dout_2[4]));
//  Memory array element: COL: 2, ROW: 5
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_101(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[5]), .O(pre_dout_2[5]));
//  Memory array element: COL: 2, ROW: 6
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_102(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[6]), .O(pre_dout_2[6]));
//  Memory array element: COL: 2, ROW: 7
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_103(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[7]), .O(pre_dout_2[7]));
//  Memory array element: COL: 2, ROW: 8
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_104(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[8]), .O(pre_dout_2[8]));
//  Memory array element: COL: 2, ROW: 9
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_105(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[9]), .O(pre_dout_2[9]));
//  Memory array element: COL: 2, ROW: 10
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_106(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[10]), .O(pre_dout_2[10]));
//  Memory array element: COL: 2, ROW: 11
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_107(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[11]), .O(pre_dout_2[11]));
//  Memory array element: COL: 2, ROW: 12
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_108(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[12]), .O(pre_dout_2[12]));
//  Memory array element: COL: 2, ROW: 13
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_109(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[13]), .O(pre_dout_2[13]));
//  Memory array element: COL: 2, ROW: 14
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_110(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[14]), .O(pre_dout_2[14]));
//  Memory array element: COL: 2, ROW: 15
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_111(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[15]), .O(pre_dout_2[15]));
//  Memory array element: COL: 3, ROW: 0
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_112(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[0]), .O(pre_dout_3[0]));
//  Memory array element: COL: 3, ROW: 1
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_113(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[1]), .O(pre_dout_3[1]));
//  Memory array element: COL: 3, ROW: 2
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_114(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[2]), .O(pre_dout_3[2]));
//  Memory array element: COL: 3, ROW: 3
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_115(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[3]), .O(pre_dout_3[3]));
//  Memory array element: COL: 3, ROW: 4
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_116(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[4]), .O(pre_dout_3[4]));
//  Memory array element: COL: 3, ROW: 5
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_117(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[5]), .O(pre_dout_3[5]));
//  Memory array element: COL: 3, ROW: 6
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_118(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[6]), .O(pre_dout_3[6]));
//  Memory array element: COL: 3, ROW: 7
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_119(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[7]), .O(pre_dout_3[7]));
//  Memory array element: COL: 3, ROW: 8
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_120(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[8]), .O(pre_dout_3[8]));
//  Memory array element: COL: 3, ROW: 9
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_121(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[9]), .O(pre_dout_3[9]));
//  Memory array element: COL: 3, ROW: 10
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_122(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[10]), .O(pre_dout_3[10]));
//  Memory array element: COL: 3, ROW: 11
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_123(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[11]), .O(pre_dout_3[11]));
//  Memory array element: COL: 3, ROW: 12
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_124(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[12]), .O(pre_dout_3[12]));
//  Memory array element: COL: 3, ROW: 13
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_125(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[13]), .O(pre_dout_3[13]));
//  Memory array element: COL: 3, ROW: 14
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_126(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[14]), .O(pre_dout_3[14]));
//  Memory array element: COL: 3, ROW: 15
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_127(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[15]), .O(pre_dout_3[15]));
endmodule



module resized_HH2_xy_structuralmemory_2116ed52_(CLK_u11, bus_3407a066_, bus_02a6eccb_, bus_404a7c0c_, bus_7ff7fda2_, bus_05f7b94c_, bus_5ba84a22_, bus_084c0cb4_, bus_749f2f87_);
input		CLK_u11;
input		bus_3407a066_;
input	[31:0]	bus_02a6eccb_;
input	[2:0]	bus_404a7c0c_;
input		bus_7ff7fda2_;
input		bus_05f7b94c_;
input	[15:0]	bus_5ba84a22_;
output	[15:0]	bus_084c0cb4_;
output		bus_749f2f87_;
wire	[15:0]	bus_70deef96_;
wire		and_4f3500db_u0;
wire		or_430a5b78_u0;
wire		not_710e9279_u0;
reg		logicalMem_45d95d5f_we_delay0_u0=1'h0;
wire		or_36d51d2a_u0;
resized_HH2_xy_forge_memory_512x16_23 resized_HH2_xy_forge_memory_512x16_23_instance0(.CLK(CLK_u11), 
  .EN(or_430a5b78_u0), .WE(bus_05f7b94c_), .ADDR(bus_02a6eccb_), .DIN(bus_5ba84a22_), 
  .DOUT(bus_70deef96_), .DONE());
assign and_4f3500db_u0=bus_7ff7fda2_&not_710e9279_u0;
assign or_430a5b78_u0=bus_7ff7fda2_|bus_05f7b94c_;
assign bus_084c0cb4_=bus_70deef96_;
assign bus_749f2f87_=or_36d51d2a_u0;
assign not_710e9279_u0=~bus_05f7b94c_;
always @(posedge CLK_u11 or posedge bus_3407a066_)
begin
if (bus_3407a066_)
logicalMem_45d95d5f_we_delay0_u0<=1'h0;
else logicalMem_45d95d5f_we_delay0_u0<=bus_05f7b94c_;
end
assign or_36d51d2a_u0=and_4f3500db_u0|logicalMem_45d95d5f_we_delay0_u0;
endmodule



module resized_HH2_xy_stateVar_Out1PortEnable(bus_6395a33f_, bus_160e9142_, bus_4d5774e5_, bus_6173af9a_, bus_2635a5e4_);
input		bus_6395a33f_;
input		bus_160e9142_;
input		bus_4d5774e5_;
input		bus_6173af9a_;
output		bus_2635a5e4_;
reg		stateVar_Out1PortEnable_u1=1'h0;
assign bus_2635a5e4_=stateVar_Out1PortEnable_u1;
always @(posedge bus_6395a33f_ or posedge bus_160e9142_)
begin
if (bus_160e9142_)
stateVar_Out1PortEnable_u1<=1'h0;
else if (bus_4d5774e5_)
stateVar_Out1PortEnable_u1<=bus_6173af9a_;
end
endmodule



module resized_HH2_xy_structuralmemory_121950d1_(CLK_u12, bus_1b9eeab7_, bus_4a6c0845_, bus_0355a864_, bus_00c34d18_, bus_200222a1_, bus_4aa3f2c6_, bus_046d1002_, bus_68a9d0f3_);
input		CLK_u12;
input		bus_1b9eeab7_;
input	[31:0]	bus_4a6c0845_;
input	[2:0]	bus_0355a864_;
input		bus_00c34d18_;
input		bus_200222a1_;
input	[15:0]	bus_4aa3f2c6_;
output	[15:0]	bus_046d1002_;
output		bus_68a9d0f3_;
wire	[15:0]	bus_6d117deb_;
wire		and_011ac791_u0;
wire		or_454206ee_u0;
wire		or_2c526a5c_u0;
wire		not_010b35df_u0;
reg		logicalMem_3c3a5c05_we_delay0_u0=1'h0;
resized_HH2_xy_forge_memory_512x16_23 resized_HH2_xy_forge_memory_512x16_23_instance1(.CLK(CLK_u12), 
  .EN(or_454206ee_u0), .WE(bus_200222a1_), .ADDR(bus_4a6c0845_), .DIN(bus_4aa3f2c6_), 
  .DOUT(bus_6d117deb_), .DONE());
assign and_011ac791_u0=bus_00c34d18_&not_010b35df_u0;
assign or_454206ee_u0=bus_00c34d18_|bus_200222a1_;
assign or_2c526a5c_u0=and_011ac791_u0|logicalMem_3c3a5c05_we_delay0_u0;
assign not_010b35df_u0=~bus_200222a1_;
assign bus_046d1002_=bus_6d117deb_;
assign bus_68a9d0f3_=or_2c526a5c_u0;
always @(posedge CLK_u12 or posedge bus_1b9eeab7_)
begin
if (bus_1b9eeab7_)
logicalMem_3c3a5c05_we_delay0_u0<=1'h0;
else logicalMem_3c3a5c05_we_delay0_u0<=bus_200222a1_;
end
endmodule



module resized_HH2_xy_endianswapper_6a3b12b8_(endianswapper_6a3b12b8_in, endianswapper_6a3b12b8_out);
input		endianswapper_6a3b12b8_in;
output		endianswapper_6a3b12b8_out;
assign endianswapper_6a3b12b8_out=endianswapper_6a3b12b8_in;
endmodule



module resized_HH2_xy_endianswapper_3c9180e4_(endianswapper_3c9180e4_in, endianswapper_3c9180e4_out);
input		endianswapper_3c9180e4_in;
output		endianswapper_3c9180e4_out;
assign endianswapper_3c9180e4_out=endianswapper_3c9180e4_in;
endmodule



module resized_HH2_xy_stateVar_fsmState_resized_HH2_xy(bus_027c1c08_, bus_1040e6d7_, bus_1c5da006_, bus_69c25494_, bus_6a6e976a_);
input		bus_027c1c08_;
input		bus_1040e6d7_;
input		bus_1c5da006_;
input		bus_69c25494_;
output		bus_6a6e976a_;
reg		stateVar_fsmState_resized_HH2_xy_u0=1'h0;
wire		endianswapper_6a3b12b8_out;
wire		endianswapper_3c9180e4_out;
always @(posedge bus_027c1c08_ or posedge bus_1040e6d7_)
begin
if (bus_1040e6d7_)
stateVar_fsmState_resized_HH2_xy_u0<=1'h0;
else if (bus_1c5da006_)
stateVar_fsmState_resized_HH2_xy_u0<=endianswapper_3c9180e4_out;
end
resized_HH2_xy_endianswapper_6a3b12b8_ resized_HH2_xy_endianswapper_6a3b12b8__1(.endianswapper_6a3b12b8_in(stateVar_fsmState_resized_HH2_xy_u0), 
  .endianswapper_6a3b12b8_out(endianswapper_6a3b12b8_out));
resized_HH2_xy_endianswapper_3c9180e4_ resized_HH2_xy_endianswapper_3c9180e4__1(.endianswapper_3c9180e4_in(bus_69c25494_), 
  .endianswapper_3c9180e4_out(endianswapper_3c9180e4_out));
assign bus_6a6e976a_=endianswapper_6a3b12b8_out;
endmodule



module resized_HH2_xy_endianswapper_5133b767_(endianswapper_5133b767_in, endianswapper_5133b767_out);
input	[15:0]	endianswapper_5133b767_in;
output	[15:0]	endianswapper_5133b767_out;
assign endianswapper_5133b767_out=endianswapper_5133b767_in;
endmodule



module resized_HH2_xy_endianswapper_2e0678b0_(endianswapper_2e0678b0_in, endianswapper_2e0678b0_out);
input	[15:0]	endianswapper_2e0678b0_in;
output	[15:0]	endianswapper_2e0678b0_out;
assign endianswapper_2e0678b0_out=endianswapper_2e0678b0_in;
endmodule



module resized_HH2_xy_stateVar_rowRepeated(bus_49b93211_, bus_0c3dac10_, bus_58b6be80_, bus_39234c02_, bus_4e9c8a8a_, bus_4cf3f116_, bus_3fd024dd_);
input		bus_49b93211_;
input		bus_0c3dac10_;
input		bus_58b6be80_;
input	[15:0]	bus_39234c02_;
input		bus_4e9c8a8a_;
input	[15:0]	bus_4cf3f116_;
output	[15:0]	bus_3fd024dd_;
wire	[15:0]	endianswapper_5133b767_out;
wire		or_33875961_u0;
wire	[15:0]	endianswapper_2e0678b0_out;
wire	[15:0]	mux_0e08add2_u0;
reg	[15:0]	stateVar_rowRepeated_u1=16'h1;
assign bus_3fd024dd_=endianswapper_5133b767_out;
resized_HH2_xy_endianswapper_5133b767_ resized_HH2_xy_endianswapper_5133b767__1(.endianswapper_5133b767_in(stateVar_rowRepeated_u1), 
  .endianswapper_5133b767_out(endianswapper_5133b767_out));
assign or_33875961_u0=bus_58b6be80_|bus_4e9c8a8a_;
resized_HH2_xy_endianswapper_2e0678b0_ resized_HH2_xy_endianswapper_2e0678b0__1(.endianswapper_2e0678b0_in(mux_0e08add2_u0), 
  .endianswapper_2e0678b0_out(endianswapper_2e0678b0_out));
assign mux_0e08add2_u0=(bus_58b6be80_)?bus_39234c02_:16'h1;
always @(posedge bus_49b93211_ or posedge bus_0c3dac10_)
begin
if (bus_0c3dac10_)
stateVar_rowRepeated_u1<=16'h1;
else if (or_33875961_u0)
stateVar_rowRepeated_u1<=endianswapper_2e0678b0_out;
end
endmodule



module resized_HH2_xy_endianswapper_0510eff3_(endianswapper_0510eff3_in, endianswapper_0510eff3_out);
input	[31:0]	endianswapper_0510eff3_in;
output	[31:0]	endianswapper_0510eff3_out;
assign endianswapper_0510eff3_out=endianswapper_0510eff3_in;
endmodule



module resized_HH2_xy_endianswapper_2b65c73c_(endianswapper_2b65c73c_in, endianswapper_2b65c73c_out);
input	[31:0]	endianswapper_2b65c73c_in;
output	[31:0]	endianswapper_2b65c73c_out;
assign endianswapper_2b65c73c_out=endianswapper_2b65c73c_in;
endmodule



module resized_HH2_xy_stateVar_Out1MaxTokenIndex(bus_2fb5cc44_, bus_2eaa1fa7_, bus_0662c425_, bus_799d8f37_, bus_0b94f26f_);
input		bus_2fb5cc44_;
input		bus_2eaa1fa7_;
input		bus_0662c425_;
input	[31:0]	bus_799d8f37_;
output	[31:0]	bus_0b94f26f_;
wire	[31:0]	endianswapper_0510eff3_out;
wire	[31:0]	endianswapper_2b65c73c_out;
reg	[31:0]	stateVar_Out1MaxTokenIndex_u1=32'h0;
assign bus_0b94f26f_=endianswapper_0510eff3_out;
resized_HH2_xy_endianswapper_0510eff3_ resized_HH2_xy_endianswapper_0510eff3__1(.endianswapper_0510eff3_in(stateVar_Out1MaxTokenIndex_u1), 
  .endianswapper_0510eff3_out(endianswapper_0510eff3_out));
resized_HH2_xy_endianswapper_2b65c73c_ resized_HH2_xy_endianswapper_2b65c73c__1(.endianswapper_2b65c73c_in(bus_799d8f37_), 
  .endianswapper_2b65c73c_out(endianswapper_2b65c73c_out));
always @(posedge bus_2fb5cc44_ or posedge bus_2eaa1fa7_)
begin
if (bus_2eaa1fa7_)
stateVar_Out1MaxTokenIndex_u1<=32'h0;
else if (bus_0662c425_)
stateVar_Out1MaxTokenIndex_u1<=endianswapper_2b65c73c_out;
end
endmodule



module resized_HH2_xy_endianswapper_1059625e_(endianswapper_1059625e_in, endianswapper_1059625e_out);
input	[15:0]	endianswapper_1059625e_in;
output	[15:0]	endianswapper_1059625e_out;
assign endianswapper_1059625e_out=endianswapper_1059625e_in;
endmodule



module resized_HH2_xy_endianswapper_4f7ac960_(endianswapper_4f7ac960_in, endianswapper_4f7ac960_out);
input	[15:0]	endianswapper_4f7ac960_in;
output	[15:0]	endianswapper_4f7ac960_out;
assign endianswapper_4f7ac960_out=endianswapper_4f7ac960_in;
endmodule



module resized_HH2_xy_stateVar_x(bus_2e51ce68_, bus_365ac0ca_, bus_5f0f6c4a_, bus_1f3118e6_, bus_2341ca1a_, bus_25e6f202_, bus_5931117b_);
input		bus_2e51ce68_;
input		bus_365ac0ca_;
input		bus_5f0f6c4a_;
input	[15:0]	bus_1f3118e6_;
input		bus_2341ca1a_;
input	[15:0]	bus_25e6f202_;
output	[15:0]	bus_5931117b_;
wire	[15:0]	mux_5f009b90_u0;
wire		or_24f369a7_u0;
reg	[15:0]	stateVar_x_u1=16'h0;
wire	[15:0]	endianswapper_1059625e_out;
wire	[15:0]	endianswapper_4f7ac960_out;
assign mux_5f009b90_u0=(bus_5f0f6c4a_)?bus_1f3118e6_:16'h0;
assign or_24f369a7_u0=bus_5f0f6c4a_|bus_2341ca1a_;
always @(posedge bus_2e51ce68_ or posedge bus_365ac0ca_)
begin
if (bus_365ac0ca_)
stateVar_x_u1<=16'h0;
else if (or_24f369a7_u0)
stateVar_x_u1<=endianswapper_1059625e_out;
end
assign bus_5931117b_=endianswapper_4f7ac960_out;
resized_HH2_xy_endianswapper_1059625e_ resized_HH2_xy_endianswapper_1059625e__1(.endianswapper_1059625e_in(mux_5f009b90_u0), 
  .endianswapper_1059625e_out(endianswapper_1059625e_out));
resized_HH2_xy_endianswapper_4f7ac960_ resized_HH2_xy_endianswapper_4f7ac960__1(.endianswapper_4f7ac960_in(stateVar_x_u1), 
  .endianswapper_4f7ac960_out(endianswapper_4f7ac960_out));
endmodule



module resized_HH2_xy_endianswapper_6888af0b_(endianswapper_6888af0b_in, endianswapper_6888af0b_out);
input	[31:0]	endianswapper_6888af0b_in;
output	[31:0]	endianswapper_6888af0b_out;
assign endianswapper_6888af0b_out=32'h0;
endmodule



module resized_HH2_xy_endianswapper_52dc6dda_(endianswapper_52dc6dda_in, endianswapper_52dc6dda_out);
input	[31:0]	endianswapper_52dc6dda_in;
output	[31:0]	endianswapper_52dc6dda_out;
assign endianswapper_52dc6dda_out=32'h0;
endmodule



module resized_HH2_xy_stateVar_fsmOldState_resized_HH2_xy(bus_5900bf5a_, bus_353bfc63_, bus_58660ccc_, bus_6ef2aeea_, bus_2ae1483e_);
input		bus_5900bf5a_;
input		bus_353bfc63_;
input		bus_58660ccc_;
input	[31:0]	bus_6ef2aeea_;
output	[31:0]	bus_2ae1483e_;
wire	[31:0]	endianswapper_6888af0b_out;
wire	[31:0]	endianswapper_52dc6dda_out;
resized_HH2_xy_endianswapper_6888af0b_ resized_HH2_xy_endianswapper_6888af0b__1(.endianswapper_6888af0b_in(32'h0), 
  .endianswapper_6888af0b_out(endianswapper_6888af0b_out));
resized_HH2_xy_endianswapper_52dc6dda_ resized_HH2_xy_endianswapper_52dc6dda__1(.endianswapper_52dc6dda_in(32'h0), 
  .endianswapper_52dc6dda_out(endianswapper_52dc6dda_out));
assign bus_2ae1483e_=32'h0;
endmodule



module resized_HH2_xy_simplememoryreferee_390f3e2f_(bus_23993a97_, bus_7cef1f98_, bus_7ebc765f_, bus_2d8c8d97_, bus_71cc810b_, bus_7a8a14d8_, bus_706609c9_, bus_2df6d93b_, bus_2ded108e_, bus_2e3a2c30_, bus_14e3e00d_, bus_194afe2d_, bus_647b7d66_, bus_4b65d917_, bus_4edd6dce_, bus_7a3d3bb9_, bus_46701177_, bus_1caadeaa_, bus_480a5dc4_, bus_43e739c0_, bus_70595e48_, bus_37b58ffd_, bus_7faadc73_, bus_6ae64912_);
input		bus_23993a97_;
input		bus_7cef1f98_;
input		bus_7ebc765f_;
input	[15:0]	bus_2d8c8d97_;
input		bus_71cc810b_;
input	[15:0]	bus_7a8a14d8_;
input	[31:0]	bus_706609c9_;
input	[2:0]	bus_2df6d93b_;
input		bus_2ded108e_;
input	[15:0]	bus_2e3a2c30_;
input	[31:0]	bus_14e3e00d_;
input	[2:0]	bus_194afe2d_;
input		bus_647b7d66_;
input	[31:0]	bus_4b65d917_;
input	[2:0]	bus_4edd6dce_;
output	[15:0]	bus_7a3d3bb9_;
output	[31:0]	bus_46701177_;
output		bus_1caadeaa_;
output		bus_480a5dc4_;
output	[2:0]	bus_43e739c0_;
output		bus_70595e48_;
output		bus_37b58ffd_;
output	[15:0]	bus_7faadc73_;
output		bus_6ae64912_;
wire	[15:0]	mux_438ddb2c_u0;
reg		done_qual_u105=1'h0;
reg		done_qual_u106_u0=1'h0;
wire		not_78100a33_u0;
wire	[31:0]	mux_2cce096b_u0;
wire		not_4368e9cf_u0;
reg		done_qual_u107_u0=1'h0;
wire		and_2ace2342_u0;
wire		and_398a441b_u0;
wire		or_6ce15fd9_u0;
wire		or_32a03c19_u0;
wire		not_60905529_u0;
wire		or_3056934c_u0;
wire		or_5f2fcc54_u0;
wire		and_3175db2e_u0;
wire		or_7c3a72c7_u0;
assign mux_438ddb2c_u0=(bus_71cc810b_)?bus_7a8a14d8_:bus_2e3a2c30_;
always @(posedge bus_23993a97_)
begin
if (bus_7cef1f98_)
done_qual_u105<=1'h0;
else done_qual_u105<=bus_647b7d66_;
end
always @(posedge bus_23993a97_)
begin
if (bus_7cef1f98_)
done_qual_u106_u0<=1'h0;
else done_qual_u106_u0<=bus_71cc810b_;
end
assign not_78100a33_u0=~bus_7ebc765f_;
assign mux_2cce096b_u0=({32{bus_71cc810b_}}&bus_706609c9_)|({32{bus_2ded108e_}}&bus_14e3e00d_)|({32{bus_647b7d66_}}&bus_4b65d917_);
assign not_4368e9cf_u0=~bus_7ebc765f_;
always @(posedge bus_23993a97_)
begin
if (bus_7cef1f98_)
done_qual_u107_u0<=1'h0;
else done_qual_u107_u0<=bus_2ded108e_;
end
assign and_2ace2342_u0=or_32a03c19_u0&bus_7ebc765f_;
assign bus_7a3d3bb9_=mux_438ddb2c_u0;
assign bus_46701177_=mux_2cce096b_u0;
assign bus_1caadeaa_=or_6ce15fd9_u0;
assign bus_480a5dc4_=or_5f2fcc54_u0;
assign bus_43e739c0_=3'h1;
assign bus_70595e48_=and_2ace2342_u0;
assign bus_37b58ffd_=and_398a441b_u0;
assign bus_7faadc73_=bus_2d8c8d97_;
assign bus_6ae64912_=and_3175db2e_u0;
assign and_398a441b_u0=or_3056934c_u0&bus_7ebc765f_;
assign or_6ce15fd9_u0=bus_71cc810b_|bus_2ded108e_;
assign or_32a03c19_u0=bus_71cc810b_|done_qual_u106_u0;
assign not_60905529_u0=~bus_7ebc765f_;
assign or_3056934c_u0=bus_2ded108e_|done_qual_u107_u0;
assign or_5f2fcc54_u0=bus_71cc810b_|bus_2ded108e_|bus_647b7d66_;
assign and_3175db2e_u0=or_7c3a72c7_u0&bus_7ebc765f_;
assign or_7c3a72c7_u0=bus_647b7d66_|done_qual_u105;
endmodule



module resized_HH2_xy_consumeRow(CLK, RESET, GO, port_0bc8ac8b_, port_3de2b1d0_, port_01480d6c_, port_43c4e7d2_, RESULT, RESULT_u1352, RESULT_u1353, RESULT_u1354, RESULT_u1355, RESULT_u1356, RESULT_u1357, RESULT_u1358, RESULT_u1359, RESULT_u1360, RESULT_u1361, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_0bc8ac8b_;
input		port_3de2b1d0_;
input		port_01480d6c_;
input	[15:0]	port_43c4e7d2_;
output		RESULT;
output	[15:0]	RESULT_u1352;
output		RESULT_u1353;
output	[31:0]	RESULT_u1354;
output	[15:0]	RESULT_u1355;
output	[2:0]	RESULT_u1356;
output		RESULT_u1357;
output	[31:0]	RESULT_u1358;
output	[15:0]	RESULT_u1359;
output	[2:0]	RESULT_u1360;
output		RESULT_u1361;
output		DONE;
wire		simplePinWrite;
wire signed	[16:0]	lessThanEqualTo_b_signed;
wire		lessThanEqualTo;
wire signed	[16:0]	lessThanEqualTo_a_signed;
wire		and_u2243_u0;
wire		and_u2244_u0;
wire		not_u413_u0;
wire	[31:0]	add;
wire	[31:0]	add_u168;
reg		reg_4491e8e1_u0=1'h0;
wire		and_u2245_u0;
wire		or_u708_u0;
wire	[15:0]	add_u169;
reg	[15:0]	syncEnable_u326=16'h0;
wire		and_u2246_u0;
wire		and_u2247_u0;
reg		and_delayed_u149=1'h0;
wire	[15:0]	mux_u244;
wire	[15:0]	latch_6c179c2e_out;
reg	[15:0]	latch_6c179c2e_reg=16'h0;
wire		or_u709_u0;
wire	[15:0]	add_u170;
wire		and_u2248_u0;
wire signed	[16:0]	lessThanEqualTo_u1_a_signed;
wire signed	[16:0]	lessThanEqualTo_u1_b_signed;
wire		lessThanEqualTo_u1;
wire		and_u2249_u0;
wire		not_u414_u0;
wire		and_u2250_u0;
reg		and_delayed_u150_u0=1'h0;
wire		and_u2251_u0;
wire	[15:0]	subtract;
wire	[31:0]	add_u171;
reg		reg_4870b88a_u0=1'h0;
wire		and_u2252_u0;
wire		or_u710_u0;
wire	[15:0]	add_u172;
reg	[15:0]	syncEnable_u327_u0=16'h0;
wire	[15:0]	latch_3f25af03_out;
reg	[15:0]	latch_3f25af03_reg=16'h0;
wire	[15:0]	mux_u245_u0;
wire		or_u711_u0;
reg	[15:0]	syncEnable_u328_u0=16'h0;
reg		reg_34ad0c93_u0=1'h0;
assign simplePinWrite=GO&{1{GO}};
assign lessThanEqualTo_a_signed={mux_u244[15], mux_u244};
assign lessThanEqualTo_b_signed=17'h3;
assign lessThanEqualTo=lessThanEqualTo_a_signed<=lessThanEqualTo_b_signed;
assign and_u2243_u0=or_u709_u0&not_u413_u0;
assign and_u2244_u0=or_u709_u0&lessThanEqualTo;
assign not_u413_u0=~lessThanEqualTo;
assign add={14'b0, port_0bc8ac8b_, 2'b0}+{mux_u244[15], mux_u244[15], mux_u244[15], mux_u244[15], mux_u244[15], mux_u244[15], mux_u244[15], mux_u244[15], mux_u244[15], mux_u244[15], mux_u244[15], mux_u244[15], mux_u244[15], mux_u244[15], mux_u244[15], mux_u244[15], mux_u244};
assign add_u168={add[19], add[19], add[19], add[19], add[19], add[19], add[19], add[19], add[19], add[19], add[19], add[19], add[19:0]}+32'h0;
always @(posedge CLK or posedge and_u2247_u0 or posedge or_u708_u0)
begin
if (or_u708_u0)
reg_4491e8e1_u0<=1'h0;
else if (and_u2247_u0)
reg_4491e8e1_u0<=1'h1;
else reg_4491e8e1_u0<=reg_4491e8e1_u0;
end
assign and_u2245_u0=reg_4491e8e1_u0&port_3de2b1d0_;
assign or_u708_u0=and_u2245_u0|RESET;
assign add_u169=mux_u244+16'h1;
always @(posedge CLK)
begin
if (and_u2247_u0)
syncEnable_u326<=add_u169;
end
assign and_u2246_u0=and_u2243_u0&or_u709_u0;
assign and_u2247_u0=and_u2244_u0&or_u709_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u149<=1'h0;
else and_delayed_u149<=and_u2247_u0;
end
assign mux_u244=(GO)?16'h0:syncEnable_u326;
assign latch_6c179c2e_out=(GO)?port_43c4e7d2_:latch_6c179c2e_reg;
always @(posedge CLK)
begin
if (GO)
latch_6c179c2e_reg<=port_43c4e7d2_;
end
assign or_u709_u0=GO|and_delayed_u149;
assign add_u170=port_0bc8ac8b_+16'h1;
assign and_u2248_u0=and_u2250_u0&or_u711_u0;
assign lessThanEqualTo_u1_a_signed={mux_u245_u0[15], mux_u245_u0};
assign lessThanEqualTo_u1_b_signed=17'h4;
assign lessThanEqualTo_u1=lessThanEqualTo_u1_a_signed<=lessThanEqualTo_u1_b_signed;
assign and_u2249_u0=or_u711_u0&not_u414_u0;
assign not_u414_u0=~lessThanEqualTo_u1;
assign and_u2250_u0=or_u711_u0&lessThanEqualTo_u1;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u150_u0<=1'h0;
else and_delayed_u150_u0<=and_u2248_u0;
end
assign and_u2251_u0=and_u2249_u0&or_u711_u0;
assign subtract=mux_u245_u0-16'h1;
assign add_u171={subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract}+32'h0;
always @(posedge CLK or posedge and_u2248_u0 or posedge or_u710_u0)
begin
if (or_u710_u0)
reg_4870b88a_u0<=1'h0;
else if (and_u2248_u0)
reg_4870b88a_u0<=1'h1;
else reg_4870b88a_u0<=reg_4870b88a_u0;
end
assign and_u2252_u0=reg_4870b88a_u0&port_01480d6c_;
assign or_u710_u0=and_u2252_u0|RESET;
assign add_u172=mux_u245_u0+16'h1;
always @(posedge CLK)
begin
if (and_u2248_u0)
syncEnable_u327_u0<=add_u172;
end
assign latch_3f25af03_out=(GO)?port_43c4e7d2_:latch_3f25af03_reg;
always @(posedge CLK)
begin
if (GO)
latch_3f25af03_reg<=port_43c4e7d2_;
end
assign mux_u245_u0=(GO)?16'h1:syncEnable_u327_u0;
assign or_u711_u0=GO|and_delayed_u150_u0;
always @(posedge CLK)
begin
if (GO)
syncEnable_u328_u0<=add_u170;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_34ad0c93_u0<=1'h0;
else reg_34ad0c93_u0<=and_u2246_u0;
end
assign RESULT=and_u2246_u0;
assign RESULT_u1352=syncEnable_u328_u0;
assign RESULT_u1353=and_u2247_u0;
assign RESULT_u1354=add_u168;
assign RESULT_u1355=latch_6c179c2e_out;
assign RESULT_u1356=3'h1;
assign RESULT_u1357=and_u2248_u0;
assign RESULT_u1358=add_u171;
assign RESULT_u1359=latch_3f25af03_out;
assign RESULT_u1360=3'h1;
assign RESULT_u1361=simplePinWrite;
assign DONE=reg_34ad0c93_u0;
endmodule



module resized_HH2_xy_repeatRowExpanded(CLK, RESET, GO, port_3ddff29c_, port_42abce2f_, port_6af401d3_, port_516974d5_, RESULT, RESULT_u1362, RESULT_u1363, RESULT_u1364, RESULT_u1365, RESULT_u1366, RESULT_u1367, RESULT_u1368, RESULT_u1369, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_3ddff29c_;
input		port_42abce2f_;
input	[15:0]	port_6af401d3_;
input		port_516974d5_;
output		RESULT;
output	[15:0]	RESULT_u1362;
output		RESULT_u1363;
output	[31:0]	RESULT_u1364;
output	[2:0]	RESULT_u1365;
output		RESULT_u1366;
output	[31:0]	RESULT_u1367;
output	[15:0]	RESULT_u1368;
output	[2:0]	RESULT_u1369;
output		DONE;
wire	[15:0]	add;
wire		and_u2253_u0;
reg		and_delayed_u151=1'h0;
wire signed	[31:0]	lessThan_b_signed;
wire signed	[31:0]	lessThan_a_signed;
wire		lessThan;
wire		and_u2254_u0;
wire		and_u2255_u0;
wire		not_u415_u0;
wire	[31:0]	add_u173;
wire		and_u2256_u0;
wire	[31:0]	add_u174;
wire		and_u2257_u0;
reg		reg_1786c6a0_u0=1'h0;
wire		or_u712_u0;
wire	[31:0]	add_u175;
reg	[31:0]	syncEnable_u329=32'h0;
wire		and_u2258_u0;
wire	[31:0]	mux_u246;
wire		or_u713_u0;
reg		reg_48f0c82f_u0=1'h0;
assign add=port_3ddff29c_+16'h1;
assign and_u2253_u0=and_u2255_u0&or_u713_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u151<=1'h0;
else and_delayed_u151<=and_u2253_u0;
end
assign lessThan_a_signed=mux_u246;
assign lessThan_b_signed=32'h200;
assign lessThan=lessThan_a_signed<lessThan_b_signed;
assign and_u2254_u0=or_u713_u0&not_u415_u0;
assign and_u2255_u0=or_u713_u0&lessThan;
assign not_u415_u0=~lessThan;
assign add_u173=mux_u246+32'h0;
assign and_u2256_u0=and_u2253_u0&port_42abce2f_;
assign add_u174=mux_u246+32'h0;
assign and_u2257_u0=reg_1786c6a0_u0&port_516974d5_;
always @(posedge CLK or posedge and_u2253_u0 or posedge or_u712_u0)
begin
if (or_u712_u0)
reg_1786c6a0_u0<=1'h0;
else if (and_u2253_u0)
reg_1786c6a0_u0<=1'h1;
else reg_1786c6a0_u0<=reg_1786c6a0_u0;
end
assign or_u712_u0=and_u2257_u0|RESET;
assign add_u175=mux_u246+32'h1;
always @(posedge CLK)
begin
if (and_u2253_u0)
syncEnable_u329<=add_u175;
end
assign and_u2258_u0=and_u2254_u0&or_u713_u0;
assign mux_u246=(reg_48f0c82f_u0)?32'h0:syncEnable_u329;
assign or_u713_u0=reg_48f0c82f_u0|and_delayed_u151;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_48f0c82f_u0<=1'h0;
else reg_48f0c82f_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u1362=add;
assign RESULT_u1363=and_u2253_u0;
assign RESULT_u1364=add_u173;
assign RESULT_u1365=3'h1;
assign RESULT_u1366=and_u2253_u0;
assign RESULT_u1367=add_u174;
assign RESULT_u1368=port_6af401d3_;
assign RESULT_u1369=3'h1;
assign DONE=and_u2258_u0;
endmodule



module resized_HH2_xy_globalreset_physical_08a74754_(bus_139efad7_, bus_67634e72_, bus_0b61c797_);
input		bus_139efad7_;
input		bus_67634e72_;
output		bus_0b61c797_;
reg		sample_u35=1'h0;
reg		cross_u35=1'h0;
reg		glitch_u35=1'h0;
wire		or_7c85da08_u0;
wire		and_734ae8f4_u0;
wire		not_66f3cc0d_u0;
reg		final_u35=1'h1;
always @(posedge bus_139efad7_)
begin
sample_u35<=1'h1;
end
assign bus_0b61c797_=or_7c85da08_u0;
always @(posedge bus_139efad7_)
begin
cross_u35<=sample_u35;
end
always @(posedge bus_139efad7_)
begin
glitch_u35<=cross_u35;
end
assign or_7c85da08_u0=bus_67634e72_|final_u35;
assign and_734ae8f4_u0=cross_u35&glitch_u35;
assign not_66f3cc0d_u0=~and_734ae8f4_u0;
always @(posedge bus_139efad7_)
begin
final_u35<=not_66f3cc0d_u0;
end
endmodule



module resized_HH2_xy_simplememoryreferee_519aba6e_(bus_31e46996_, bus_78041c94_, bus_69efc929_, bus_09bbc993_, bus_3ec76267_, bus_4f50e209_, bus_3cbefa4e_, bus_57eee443_, bus_5133aa26_, bus_649a3ec9_, bus_7184d705_, bus_27c6803d_, bus_5fed9ad9_, bus_1b9989aa_, bus_2570462b_, bus_13e0228b_, bus_15d988f3_, bus_08f43ee3_, bus_7fa5bd8d_);
input		bus_31e46996_;
input		bus_78041c94_;
input		bus_69efc929_;
input	[15:0]	bus_09bbc993_;
input		bus_3ec76267_;
input	[15:0]	bus_4f50e209_;
input	[31:0]	bus_3cbefa4e_;
input	[2:0]	bus_57eee443_;
input		bus_5133aa26_;
input	[31:0]	bus_649a3ec9_;
input	[2:0]	bus_7184d705_;
output	[15:0]	bus_27c6803d_;
output	[31:0]	bus_5fed9ad9_;
output		bus_1b9989aa_;
output		bus_2570462b_;
output	[2:0]	bus_13e0228b_;
output		bus_15d988f3_;
output	[15:0]	bus_08f43ee3_;
output		bus_7fa5bd8d_;
wire	[31:0]	mux_541091d0_u0;
wire		or_3c8a910a_u0;
wire		and_73495169_u0;
wire	[15:0]	mux_07bd52f9_u0;
wire		not_7c11c578_u0;
reg		done_qual_u108_u0=1'h0;
wire		not_621ffbb4_u0;
wire		and_6ff00e7d_u0;
wire		or_5eeb369c_u0;
reg		done_qual_u109_u0=1'h0;
wire		or_26f3a929_u0;
assign mux_541091d0_u0=(bus_3ec76267_)?bus_3cbefa4e_:bus_649a3ec9_;
assign or_3c8a910a_u0=bus_3ec76267_|bus_5133aa26_;
assign and_73495169_u0=or_5eeb369c_u0&bus_69efc929_;
assign mux_07bd52f9_u0=({16{bus_3ec76267_}}&bus_4f50e209_);
assign not_7c11c578_u0=~bus_69efc929_;
always @(posedge bus_31e46996_)
begin
if (bus_78041c94_)
done_qual_u108_u0<=1'h0;
else done_qual_u108_u0<=bus_3ec76267_;
end
assign not_621ffbb4_u0=~bus_69efc929_;
assign and_6ff00e7d_u0=or_26f3a929_u0&bus_69efc929_;
assign or_5eeb369c_u0=bus_5133aa26_|done_qual_u109_u0;
always @(posedge bus_31e46996_)
begin
if (bus_78041c94_)
done_qual_u109_u0<=1'h0;
else done_qual_u109_u0<=bus_5133aa26_;
end
assign or_26f3a929_u0=bus_3ec76267_|done_qual_u108_u0;
assign bus_27c6803d_=mux_07bd52f9_u0;
assign bus_5fed9ad9_=mux_541091d0_u0;
assign bus_1b9989aa_=bus_3ec76267_;
assign bus_2570462b_=or_3c8a910a_u0;
assign bus_13e0228b_=3'h1;
assign bus_15d988f3_=and_6ff00e7d_u0;
assign bus_08f43ee3_=bus_09bbc993_;
assign bus_7fa5bd8d_=and_73495169_u0;
endmodule



module resized_HH2_xy_reset(CLK, RESET, GO, RESULT, RESULT_u1370, RESULT_u1371, RESULT_u1372, DONE);
input		CLK;
input		RESET;
input		GO;
output		RESULT;
output	[15:0]	RESULT_u1370;
output		RESULT_u1371;
output	[15:0]	RESULT_u1372;
output		DONE;
reg		reg_08fe6a7b_u0=1'h0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_08fe6a7b_u0<=1'h0;
else reg_08fe6a7b_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u1370=16'h1;
assign RESULT_u1371=GO;
assign RESULT_u1372=16'h0;
assign DONE=reg_08fe6a7b_u0;
endmodule


