// __  ___ __ ___  _ __   ___  ___ 
// \ \/ / '__/ _ \| '_ \ / _ \/ __|
//  >  <| | | (_) | | | | (_) \__ \
// /_/\_\_|  \___/|_| |_|\___/|___/
// 
// Xronos synthesizer version
// Run date: Thu 2 Nov 2017 13:59:05 +0000
// 

module resized_HH3_xy(CLK, In1_ACK, In1_SEND, Out1_SEND, In1_COUNT, Out1_ACK, RESET, Out1_RDY, Out1_COUNT, Out1_DATA, In1_DATA);
wire		reset_done;
input		CLK;
output		In1_ACK;
wire		repeatRowExpanded_done;
input		In1_SEND;
wire		reset_go;
output		Out1_SEND;
input	[15:0]	In1_COUNT;
input		Out1_ACK;
wire		consumeRow_done;
input		RESET;
input		Out1_RDY;
output	[15:0]	Out1_COUNT;
wire		consumeRow_go;
output	[15:0]	Out1_DATA;
wire		repeatRowExpanded_go;
input	[15:0]	In1_DATA;
wire		bus_67ab127b_;
wire		bus_6f241b85_;
wire	[15:0]	bus_01afcb9f_;
wire		bus_368ccdf1_;
wire		reset;
wire		resized_HH3_xy_reset_instance_DONE;
wire	[15:0]	reset_u6;
wire		reset_u7;
wire	[15:0]	reset_u8;
wire		bus_402c7489_;
wire		bus_2f4398a5_;
wire	[15:0]	bus_141e2cb9_;
wire	[31:0]	bus_62beb692_;
wire		bus_461cf331_;
wire	[15:0]	bus_7b37a050_;
wire	[2:0]	bus_5740abcd_;
wire		bus_43715c56_;
wire		bus_4cfcaed6_;
wire		bus_6878fc86_;
wire		bus_0fded023_;
wire	[31:0]	bus_54879690_;
wire		bus_39aac355_;
wire	[31:0]	bus_28bc5e54_;
wire		bus_4775846d_;
wire	[15:0]	bus_27d1116c_;
wire		bus_7ca17cbb_;
wire		bus_534cc528_;
wire		bus_1a7956cb_;
wire	[2:0]	bus_55d21a89_;
wire	[15:0]	bus_0f2a4aab_;
wire		bus_75e7dd97_;
wire	[15:0]	repeatRowExpanded_u19;
wire	[2:0]	repeatRowExpanded_u20;
wire		repeatRowExpanded_u21;
wire		repeatRowExpanded;
wire		resized_HH3_xy_repeatRowExpanded_instance_DONE;
wire	[31:0]	repeatRowExpanded_u22;
wire	[2:0]	repeatRowExpanded_u23;
wire		repeatRowExpanded_u17;
wire	[31:0]	repeatRowExpanded_u18;
wire	[15:0]	repeatRowExpanded_u16;
wire	[15:0]	bus_429824b9_;
wire		bus_5fbc036a_;
wire	[15:0]	bus_1b8c04d2_;
wire		scheduler_u247;
wire		scheduler_u245;
wire	[31:0]	scheduler_u233;
wire		scheduler_u238;
wire		scheduler_u250;
wire	[31:0]	scheduler_u243;
wire		resized_HH3_xy_scheduler_instance_DONE;
wire		scheduler_u235;
wire		scheduler_u241;
wire		scheduler;
wire		scheduler_u242;
wire		scheduler_u240;
wire	[15:0]	scheduler_u249;
wire		scheduler_u236;
wire	[2:0]	scheduler_u244;
wire		scheduler_u234;
wire	[31:0]	scheduler_u239;
wire		scheduler_u248;
wire	[15:0]	scheduler_u246;
wire	[31:0]	scheduler_u237;
wire	[31:0]	bus_02dad7ef_;
wire	[31:0]	bus_6ec88e4d_;
wire	[31:0]	consumeRow_u22;
wire	[31:0]	consumeRow_u26;
wire	[2:0]	consumeRow_u28;
wire		consumeRow;
wire		consumeRow_u21;
wire	[15:0]	consumeRow_u23;
wire	[2:0]	consumeRow_u24;
wire	[15:0]	consumeRow_u27;
wire	[15:0]	consumeRow_u20;
wire		consumeRow_u25;
wire		resized_HH3_xy_consumeRow_instance_DONE;
wire		consumeRow_u29;
wire	[15:0]	bus_035cdb42_;
wire		bus_1dbe1e5d_;
assign reset_done=bus_6878fc86_;
assign In1_ACK=consumeRow_u29;
assign repeatRowExpanded_done=bus_39aac355_;
assign reset_go=scheduler_u247;
assign Out1_SEND=scheduler_u245;
assign consumeRow_done=bus_0fded023_;
assign Out1_COUNT=scheduler_u246;
assign consumeRow_go=scheduler_u248;
assign Out1_DATA=scheduler_u249;
assign repeatRowExpanded_go=scheduler_u250;
resized_HH3_xy_globalreset_physical_06d0e694_ resized_HH3_xy_globalreset_physical_06d0e694__1(.bus_647dab1e_(CLK), 
  .bus_0869a83b_(RESET), .bus_67ab127b_(bus_67ab127b_));
resized_HH3_xy_Kicker_41 resized_HH3_xy_Kicker_41_1(.CLK(CLK), .RESET(bus_67ab127b_), 
  .bus_6f241b85_(bus_6f241b85_));
resized_HH3_xy_structuralmemory_56ef0725_ resized_HH3_xy_structuralmemory_56ef0725__1(.CLK_u14(CLK), 
  .bus_5233359a_(bus_67ab127b_), .bus_4db2cf4a_(bus_62beb692_), .bus_7d712f31_(3'h1), 
  .bus_2286f07f_(bus_461cf331_), .bus_34c65aab_(bus_4cfcaed6_), .bus_25d6634e_(bus_141e2cb9_), 
  .bus_01afcb9f_(bus_01afcb9f_), .bus_368ccdf1_(bus_368ccdf1_));
resized_HH3_xy_reset resized_HH3_xy_reset_instance(.CLK(CLK), .RESET(bus_67ab127b_), 
  .GO(reset_go), .DONE(resized_HH3_xy_reset_instance_DONE), .RESULT(reset), .RESULT_u1593(reset_u6), 
  .RESULT_u1594(reset_u7), .RESULT_u1595(reset_u8));
resized_HH3_xy_simplememoryreferee_1ae795b5_ resized_HH3_xy_simplememoryreferee_1ae795b5__1(.bus_7903d426_(CLK), 
  .bus_762e0ccd_(bus_67ab127b_), .bus_12a00bf7_(bus_368ccdf1_), .bus_0d18c1eb_(bus_01afcb9f_), 
  .bus_4e950722_(consumeRow_u25), .bus_0f7eec10_(consumeRow_u27), .bus_7ccb383c_(consumeRow_u26), 
  .bus_563925df_(3'h1), .bus_2e13b093_(repeatRowExpanded_u17), .bus_75309ed5_(repeatRowExpanded_u19), 
  .bus_2c80aee2_(repeatRowExpanded_u18), .bus_104d416b_(3'h1), .bus_48029f45_(scheduler_u242), 
  .bus_0b8f5236_(scheduler_u243), .bus_4cecc8f5_(3'h1), .bus_141e2cb9_(bus_141e2cb9_), 
  .bus_62beb692_(bus_62beb692_), .bus_4cfcaed6_(bus_4cfcaed6_), .bus_461cf331_(bus_461cf331_), 
  .bus_5740abcd_(bus_5740abcd_), .bus_402c7489_(bus_402c7489_), .bus_2f4398a5_(bus_2f4398a5_), 
  .bus_7b37a050_(bus_7b37a050_), .bus_43715c56_(bus_43715c56_));
assign bus_6878fc86_=resized_HH3_xy_reset_instance_DONE&{1{resized_HH3_xy_reset_instance_DONE}};
assign bus_0fded023_=resized_HH3_xy_consumeRow_instance_DONE&{1{resized_HH3_xy_consumeRow_instance_DONE}};
resized_HH3_xy_stateVar_Out1TokenIndex resized_HH3_xy_stateVar_Out1TokenIndex_1(.bus_1a06ee5a_(CLK), 
  .bus_21fbc7d7_(bus_67ab127b_), .bus_11445d5e_(scheduler_u236), .bus_43a7b829_(scheduler_u237), 
  .bus_54879690_(bus_54879690_));
assign bus_39aac355_=resized_HH3_xy_repeatRowExpanded_instance_DONE&{1{resized_HH3_xy_repeatRowExpanded_instance_DONE}};
resized_HH3_xy_simplememoryreferee_233a65d9_ resized_HH3_xy_simplememoryreferee_233a65d9__1(.bus_0e63ff2e_(CLK), 
  .bus_2cbe6427_(bus_67ab127b_), .bus_0b7a09f9_(bus_1dbe1e5d_), .bus_3f845529_(bus_035cdb42_), 
  .bus_51dc5427_(consumeRow_u21), .bus_31d29381_(consumeRow_u23), .bus_1539b851_(consumeRow_u22), 
  .bus_5cf79b2a_(3'h1), .bus_6417eca8_(repeatRowExpanded_u21), .bus_351c3c2f_(repeatRowExpanded_u22), 
  .bus_3d2a2664_(3'h1), .bus_27d1116c_(bus_27d1116c_), .bus_28bc5e54_(bus_28bc5e54_), 
  .bus_1a7956cb_(bus_1a7956cb_), .bus_534cc528_(bus_534cc528_), .bus_55d21a89_(bus_55d21a89_), 
  .bus_4775846d_(bus_4775846d_), .bus_0f2a4aab_(bus_0f2a4aab_), .bus_7ca17cbb_(bus_7ca17cbb_));
resized_HH3_xy_stateVar_Out1PortEnable resized_HH3_xy_stateVar_Out1PortEnable_1(.bus_4966e2b3_(CLK), 
  .bus_160bb6e7_(bus_67ab127b_), .bus_4ad9d6ae_(scheduler_u240), .bus_7fa3f2df_(scheduler_u241), 
  .bus_75e7dd97_(bus_75e7dd97_));
resized_HH3_xy_repeatRowExpanded resized_HH3_xy_repeatRowExpanded_instance(.CLK(CLK), 
  .RESET(bus_67ab127b_), .GO(repeatRowExpanded_go), .port_1a399e92_(bus_1b8c04d2_), 
  .port_5a868a9f_(bus_2f4398a5_), .port_5bdc04de_(bus_7ca17cbb_), .port_095c79c5_(bus_0f2a4aab_), 
  .DONE(resized_HH3_xy_repeatRowExpanded_instance_DONE), .RESULT(repeatRowExpanded), 
  .RESULT_u1596(repeatRowExpanded_u16), .RESULT_u1600(repeatRowExpanded_u17), 
  .RESULT_u1601(repeatRowExpanded_u18), .RESULT_u1602(repeatRowExpanded_u19), 
  .RESULT_u1603(repeatRowExpanded_u20), .RESULT_u1597(repeatRowExpanded_u21), 
  .RESULT_u1598(repeatRowExpanded_u22), .RESULT_u1599(repeatRowExpanded_u23));
resized_HH3_xy_stateVar_x resized_HH3_xy_stateVar_x_1(.bus_1f8eca8a_(CLK), .bus_57b1029e_(bus_67ab127b_), 
  .bus_0ffcb094_(consumeRow), .bus_3935aade_(consumeRow_u20), .bus_1fbb8f18_(reset_u7), 
  .bus_121158f5_(16'h0), .bus_429824b9_(bus_429824b9_));
resized_HH3_xy_stateVar_fsmState_resized_HH3_xy resized_HH3_xy_stateVar_fsmState_resized_HH3_xy_1(.bus_49fba71e_(CLK), 
  .bus_1273375e_(bus_67ab127b_), .bus_0954f839_(scheduler_u234), .bus_16417063_(scheduler_u235), 
  .bus_5fbc036a_(bus_5fbc036a_));
resized_HH3_xy_stateVar_rowRepeated resized_HH3_xy_stateVar_rowRepeated_1(.bus_003a3253_(CLK), 
  .bus_7eeb9fab_(bus_67ab127b_), .bus_0e31d817_(repeatRowExpanded), .bus_7d7c11ad_(repeatRowExpanded_u16), 
  .bus_67f23a28_(reset), .bus_63962b7e_(16'h1), .bus_1b8c04d2_(bus_1b8c04d2_));
resized_HH3_xy_scheduler resized_HH3_xy_scheduler_instance(.CLK(CLK), .RESET(bus_67ab127b_), 
  .GO(bus_6f241b85_), .port_69930ca0_(32'h0), .port_7545a1a4_(bus_5fbc036a_), .port_1121f1ff_(bus_54879690_), 
  .port_70929f20_(bus_6ec88e4d_), .port_05f8f754_(bus_75e7dd97_), .port_697394d7_(bus_429824b9_), 
  .port_2ef7caed_(bus_1b8c04d2_), .port_1f63f705_(bus_43715c56_), .port_0a0e1767_(bus_7b37a050_), 
  .port_5286b1a6_(Out1_RDY), .port_64176099_(repeatRowExpanded_done), .port_21602b46_(In1_SEND), 
  .port_3915346e_(consumeRow_done), .port_3a6df956_(reset_done), .DONE(resized_HH3_xy_scheduler_instance_DONE), 
  .RESULT(scheduler), .RESULT_u1604(scheduler_u233), .RESULT_u1605(scheduler_u234), 
  .RESULT_u1606(scheduler_u235), .RESULT_u1607(scheduler_u236), .RESULT_u1608(scheduler_u237), 
  .RESULT_u1609(scheduler_u238), .RESULT_u1610(scheduler_u239), .RESULT_u1611(scheduler_u240), 
  .RESULT_u1612(scheduler_u241), .RESULT_u1613(scheduler_u242), .RESULT_u1614(scheduler_u243), 
  .RESULT_u1615(scheduler_u244), .RESULT_u1616(scheduler_u245), .RESULT_u1617(scheduler_u246), 
  .RESULT_u1618(scheduler_u247), .RESULT_u1619(scheduler_u248), .RESULT_u1620(scheduler_u249), 
  .RESULT_u1621(scheduler_u250));
resized_HH3_xy_stateVar_fsmOldState_resized_HH3_xy resized_HH3_xy_stateVar_fsmOldState_resized_HH3_xy_1(.bus_265f821d_(CLK), 
  .bus_15b24ce3_(bus_67ab127b_), .bus_4cadd642_(scheduler), .bus_11ea79c0_(32'h0), 
  .bus_02dad7ef_(bus_02dad7ef_));
resized_HH3_xy_stateVar_Out1MaxTokenIndex resized_HH3_xy_stateVar_Out1MaxTokenIndex_1(.bus_24944e90_(CLK), 
  .bus_67a2773e_(bus_67ab127b_), .bus_4329e6b2_(scheduler_u238), .bus_31a05489_(scheduler_u239), 
  .bus_6ec88e4d_(bus_6ec88e4d_));
resized_HH3_xy_consumeRow resized_HH3_xy_consumeRow_instance(.CLK(CLK), .RESET(bus_67ab127b_), 
  .GO(consumeRow_go), .port_36ed5a59_(bus_429824b9_), .port_55b6d605_(bus_4775846d_), 
  .port_7a6b4a4c_(bus_402c7489_), .port_6b0ac5ca_(In1_DATA), .DONE(resized_HH3_xy_consumeRow_instance_DONE), 
  .RESULT(consumeRow), .RESULT_u1622(consumeRow_u20), .RESULT_u1623(consumeRow_u21), 
  .RESULT_u1624(consumeRow_u22), .RESULT_u1625(consumeRow_u23), .RESULT_u1626(consumeRow_u24), 
  .RESULT_u1627(consumeRow_u25), .RESULT_u1628(consumeRow_u26), .RESULT_u1629(consumeRow_u27), 
  .RESULT_u1630(consumeRow_u28), .RESULT_u1631(consumeRow_u29));
resized_HH3_xy_structuralmemory_068f5fb6_ resized_HH3_xy_structuralmemory_068f5fb6__1(.CLK_u15(CLK), 
  .bus_13f3e3d1_(bus_67ab127b_), .bus_750d9e9a_(bus_28bc5e54_), .bus_0cd70fa4_(3'h1), 
  .bus_30fff37e_(bus_534cc528_), .bus_2ba929a7_(bus_1a7956cb_), .bus_6b58816e_(bus_27d1116c_), 
  .bus_035cdb42_(bus_035cdb42_), .bus_1dbe1e5d_(bus_1dbe1e5d_));
endmodule



module resized_HH3_xy_globalreset_physical_06d0e694_(bus_647dab1e_, bus_0869a83b_, bus_67ab127b_);
input		bus_647dab1e_;
input		bus_0869a83b_;
output		bus_67ab127b_;
reg		glitch_u37=1'h0;
reg		cross_u37=1'h0;
reg		final_u37=1'h1;
wire		or_0a2a5eff_u0;
wire		and_5ab50062_u0;
reg		sample_u37=1'h0;
wire		not_4a285c45_u0;
always @(posedge bus_647dab1e_)
begin
glitch_u37<=cross_u37;
end
always @(posedge bus_647dab1e_)
begin
cross_u37<=sample_u37;
end
always @(posedge bus_647dab1e_)
begin
final_u37<=not_4a285c45_u0;
end
assign or_0a2a5eff_u0=bus_0869a83b_|final_u37;
assign bus_67ab127b_=or_0a2a5eff_u0;
assign and_5ab50062_u0=cross_u37&glitch_u37;
always @(posedge bus_647dab1e_)
begin
sample_u37<=1'h1;
end
assign not_4a285c45_u0=~and_5ab50062_u0;
endmodule



module resized_HH3_xy_Kicker_41(CLK, RESET, bus_6f241b85_);
input		CLK;
input		RESET;
output		bus_6f241b85_;
wire		bus_19c99eae_;
wire		bus_334f4047_;
reg		kicker_2=1'h0;
wire		bus_7f3e0ffa_;
wire		bus_43a4a053_;
reg		kicker_res=1'h0;
reg		kicker_1=1'h0;
assign bus_19c99eae_=kicker_1&bus_7f3e0ffa_&bus_43a4a053_;
assign bus_334f4047_=bus_7f3e0ffa_&kicker_1;
always @(posedge CLK)
begin
kicker_2<=bus_334f4047_;
end
assign bus_7f3e0ffa_=~RESET;
assign bus_43a4a053_=~kicker_2;
always @(posedge CLK)
begin
kicker_res<=bus_19c99eae_;
end
assign bus_6f241b85_=kicker_res;
always @(posedge CLK)
begin
kicker_1<=bus_7f3e0ffa_;
end
endmodule



module resized_HH3_xy_forge_memory_512x16_28(CLK, EN, WE, ADDR, DIN, DOUT, DONE);
input		CLK;
input		EN;
input		WE;
input	[31:0]	ADDR;
input	[15:0]	DIN;
output	[15:0]	DOUT;
output		DONE;
wire		we_0;
wire	[15:0]	pre_dout_0;
wire		we_1;
wire	[15:0]	pre_dout_1;
wire		we_2;
wire	[15:0]	pre_dout_2;
wire		we_3;
wire	[15:0]	pre_dout_3;
reg	[15:0]	mux_out;
reg		wen_done;
assign we_0=WE&(ADDR[31:7]==25'h0);
assign we_1=WE&(ADDR[31:7]==25'h1);
assign we_2=WE&(ADDR[31:7]==25'h2);
assign we_3=WE&(ADDR[31:7]==25'h3);
always @(ADDR or pre_dout_0 or pre_dout_1 or pre_dout_2 or pre_dout_3)
begin
case (ADDR[31:7])25'd0:mux_out=pre_dout_0;
25'd1:mux_out=pre_dout_1;
25'd2:mux_out=pre_dout_2;
25'd3:mux_out=pre_dout_3;
default:mux_out=16'h0;
endcase end
always @(posedge CLK)
begin
wen_done<=WE;
end
assign DOUT=mux_out;
assign DONE=EN&!WE|wen_done;
//  Memory array element: COL: 0, ROW: 0
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_128(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[0]), .O(pre_dout_0[0]));
//  Memory array element: COL: 0, ROW: 1
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_129(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[1]), .O(pre_dout_0[1]));
//  Memory array element: COL: 0, ROW: 2
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_130(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[2]), .O(pre_dout_0[2]));
//  Memory array element: COL: 0, ROW: 3
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_131(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[3]), .O(pre_dout_0[3]));
//  Memory array element: COL: 0, ROW: 4
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_132(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[4]), .O(pre_dout_0[4]));
//  Memory array element: COL: 0, ROW: 5
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_133(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[5]), .O(pre_dout_0[5]));
//  Memory array element: COL: 0, ROW: 6
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_134(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[6]), .O(pre_dout_0[6]));
//  Memory array element: COL: 0, ROW: 7
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_135(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[7]), .O(pre_dout_0[7]));
//  Memory array element: COL: 0, ROW: 8
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_136(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[8]), .O(pre_dout_0[8]));
//  Memory array element: COL: 0, ROW: 9
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_137(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[9]), .O(pre_dout_0[9]));
//  Memory array element: COL: 0, ROW: 10
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_138(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[10]), .O(pre_dout_0[10]));
//  Memory array element: COL: 0, ROW: 11
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_139(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[11]), .O(pre_dout_0[11]));
//  Memory array element: COL: 0, ROW: 12
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_140(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[12]), .O(pre_dout_0[12]));
//  Memory array element: COL: 0, ROW: 13
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_141(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[13]), .O(pre_dout_0[13]));
//  Memory array element: COL: 0, ROW: 14
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_142(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[14]), .O(pre_dout_0[14]));
//  Memory array element: COL: 0, ROW: 15
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_143(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[15]), .O(pre_dout_0[15]));
//  Memory array element: COL: 1, ROW: 0
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_144(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[0]), .O(pre_dout_1[0]));
//  Memory array element: COL: 1, ROW: 1
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_145(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[1]), .O(pre_dout_1[1]));
//  Memory array element: COL: 1, ROW: 2
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_146(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[2]), .O(pre_dout_1[2]));
//  Memory array element: COL: 1, ROW: 3
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_147(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[3]), .O(pre_dout_1[3]));
//  Memory array element: COL: 1, ROW: 4
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_148(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[4]), .O(pre_dout_1[4]));
//  Memory array element: COL: 1, ROW: 5
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_149(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[5]), .O(pre_dout_1[5]));
//  Memory array element: COL: 1, ROW: 6
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_150(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[6]), .O(pre_dout_1[6]));
//  Memory array element: COL: 1, ROW: 7
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_151(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[7]), .O(pre_dout_1[7]));
//  Memory array element: COL: 1, ROW: 8
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_152(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[8]), .O(pre_dout_1[8]));
//  Memory array element: COL: 1, ROW: 9
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_153(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[9]), .O(pre_dout_1[9]));
//  Memory array element: COL: 1, ROW: 10
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_154(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[10]), .O(pre_dout_1[10]));
//  Memory array element: COL: 1, ROW: 11
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_155(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[11]), .O(pre_dout_1[11]));
//  Memory array element: COL: 1, ROW: 12
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_156(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[12]), .O(pre_dout_1[12]));
//  Memory array element: COL: 1, ROW: 13
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_157(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[13]), .O(pre_dout_1[13]));
//  Memory array element: COL: 1, ROW: 14
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_158(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[14]), .O(pre_dout_1[14]));
//  Memory array element: COL: 1, ROW: 15
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_159(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[15]), .O(pre_dout_1[15]));
//  Memory array element: COL: 2, ROW: 0
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_160(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[0]), .O(pre_dout_2[0]));
//  Memory array element: COL: 2, ROW: 1
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_161(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[1]), .O(pre_dout_2[1]));
//  Memory array element: COL: 2, ROW: 2
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_162(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[2]), .O(pre_dout_2[2]));
//  Memory array element: COL: 2, ROW: 3
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_163(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[3]), .O(pre_dout_2[3]));
//  Memory array element: COL: 2, ROW: 4
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_164(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[4]), .O(pre_dout_2[4]));
//  Memory array element: COL: 2, ROW: 5
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_165(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[5]), .O(pre_dout_2[5]));
//  Memory array element: COL: 2, ROW: 6
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_166(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[6]), .O(pre_dout_2[6]));
//  Memory array element: COL: 2, ROW: 7
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_167(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[7]), .O(pre_dout_2[7]));
//  Memory array element: COL: 2, ROW: 8
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_168(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[8]), .O(pre_dout_2[8]));
//  Memory array element: COL: 2, ROW: 9
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_169(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[9]), .O(pre_dout_2[9]));
//  Memory array element: COL: 2, ROW: 10
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_170(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[10]), .O(pre_dout_2[10]));
//  Memory array element: COL: 2, ROW: 11
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_171(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[11]), .O(pre_dout_2[11]));
//  Memory array element: COL: 2, ROW: 12
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_172(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[12]), .O(pre_dout_2[12]));
//  Memory array element: COL: 2, ROW: 13
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_173(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[13]), .O(pre_dout_2[13]));
//  Memory array element: COL: 2, ROW: 14
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_174(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[14]), .O(pre_dout_2[14]));
//  Memory array element: COL: 2, ROW: 15
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_175(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[15]), .O(pre_dout_2[15]));
//  Memory array element: COL: 3, ROW: 0
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_176(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[0]), .O(pre_dout_3[0]));
//  Memory array element: COL: 3, ROW: 1
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_177(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[1]), .O(pre_dout_3[1]));
//  Memory array element: COL: 3, ROW: 2
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_178(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[2]), .O(pre_dout_3[2]));
//  Memory array element: COL: 3, ROW: 3
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_179(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[3]), .O(pre_dout_3[3]));
//  Memory array element: COL: 3, ROW: 4
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_180(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[4]), .O(pre_dout_3[4]));
//  Memory array element: COL: 3, ROW: 5
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_181(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[5]), .O(pre_dout_3[5]));
//  Memory array element: COL: 3, ROW: 6
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_182(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[6]), .O(pre_dout_3[6]));
//  Memory array element: COL: 3, ROW: 7
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_183(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[7]), .O(pre_dout_3[7]));
//  Memory array element: COL: 3, ROW: 8
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_184(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[8]), .O(pre_dout_3[8]));
//  Memory array element: COL: 3, ROW: 9
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_185(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[9]), .O(pre_dout_3[9]));
//  Memory array element: COL: 3, ROW: 10
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_186(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[10]), .O(pre_dout_3[10]));
//  Memory array element: COL: 3, ROW: 11
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_187(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[11]), .O(pre_dout_3[11]));
//  Memory array element: COL: 3, ROW: 12
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_188(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[12]), .O(pre_dout_3[12]));
//  Memory array element: COL: 3, ROW: 13
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_189(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[13]), .O(pre_dout_3[13]));
//  Memory array element: COL: 3, ROW: 14
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_190(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[14]), .O(pre_dout_3[14]));
//  Memory array element: COL: 3, ROW: 15
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_191(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[15]), .O(pre_dout_3[15]));
endmodule



module resized_HH3_xy_structuralmemory_56ef0725_(CLK_u14, bus_5233359a_, bus_4db2cf4a_, bus_7d712f31_, bus_2286f07f_, bus_34c65aab_, bus_25d6634e_, bus_01afcb9f_, bus_368ccdf1_);
input		CLK_u14;
input		bus_5233359a_;
input	[31:0]	bus_4db2cf4a_;
input	[2:0]	bus_7d712f31_;
input		bus_2286f07f_;
input		bus_34c65aab_;
input	[15:0]	bus_25d6634e_;
output	[15:0]	bus_01afcb9f_;
output		bus_368ccdf1_;
wire		not_77c7b903_u0;
reg		logicalMem_85a5964_we_delay0_u0=1'h0;
wire	[15:0]	bus_68f904c0_;
wire		and_3328c033_u0;
wire		or_7652062c_u0;
wire		or_00a5a73a_u0;
assign not_77c7b903_u0=~bus_34c65aab_;
always @(posedge CLK_u14 or posedge bus_5233359a_)
begin
if (bus_5233359a_)
logicalMem_85a5964_we_delay0_u0<=1'h0;
else logicalMem_85a5964_we_delay0_u0<=bus_34c65aab_;
end
resized_HH3_xy_forge_memory_512x16_28 resized_HH3_xy_forge_memory_512x16_28_instance0(.CLK(CLK_u14), 
  .EN(or_00a5a73a_u0), .WE(bus_34c65aab_), .ADDR(bus_4db2cf4a_), .DIN(bus_25d6634e_), 
  .DOUT(bus_68f904c0_), .DONE());
assign bus_01afcb9f_=bus_68f904c0_;
assign bus_368ccdf1_=or_7652062c_u0;
assign and_3328c033_u0=bus_2286f07f_&not_77c7b903_u0;
assign or_7652062c_u0=and_3328c033_u0|logicalMem_85a5964_we_delay0_u0;
assign or_00a5a73a_u0=bus_2286f07f_|bus_34c65aab_;
endmodule



module resized_HH3_xy_reset(CLK, RESET, GO, RESULT, RESULT_u1593, RESULT_u1594, RESULT_u1595, DONE);
input		CLK;
input		RESET;
input		GO;
output		RESULT;
output	[15:0]	RESULT_u1593;
output		RESULT_u1594;
output	[15:0]	RESULT_u1595;
output		DONE;
reg		reg_33a87f54_u0=1'h0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_33a87f54_u0<=1'h0;
else reg_33a87f54_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u1593=16'h1;
assign RESULT_u1594=GO;
assign RESULT_u1595=16'h0;
assign DONE=reg_33a87f54_u0;
endmodule



module resized_HH3_xy_simplememoryreferee_1ae795b5_(bus_7903d426_, bus_762e0ccd_, bus_12a00bf7_, bus_0d18c1eb_, bus_4e950722_, bus_0f7eec10_, bus_7ccb383c_, bus_563925df_, bus_2e13b093_, bus_75309ed5_, bus_2c80aee2_, bus_104d416b_, bus_48029f45_, bus_0b8f5236_, bus_4cecc8f5_, bus_141e2cb9_, bus_62beb692_, bus_4cfcaed6_, bus_461cf331_, bus_5740abcd_, bus_402c7489_, bus_2f4398a5_, bus_7b37a050_, bus_43715c56_);
input		bus_7903d426_;
input		bus_762e0ccd_;
input		bus_12a00bf7_;
input	[15:0]	bus_0d18c1eb_;
input		bus_4e950722_;
input	[15:0]	bus_0f7eec10_;
input	[31:0]	bus_7ccb383c_;
input	[2:0]	bus_563925df_;
input		bus_2e13b093_;
input	[15:0]	bus_75309ed5_;
input	[31:0]	bus_2c80aee2_;
input	[2:0]	bus_104d416b_;
input		bus_48029f45_;
input	[31:0]	bus_0b8f5236_;
input	[2:0]	bus_4cecc8f5_;
output	[15:0]	bus_141e2cb9_;
output	[31:0]	bus_62beb692_;
output		bus_4cfcaed6_;
output		bus_461cf331_;
output	[2:0]	bus_5740abcd_;
output		bus_402c7489_;
output		bus_2f4398a5_;
output	[15:0]	bus_7b37a050_;
output		bus_43715c56_;
wire		and_58fc57bc_u0;
wire		or_61208902_u0;
wire		or_6978c77b_u0;
wire		or_66105f34_u0;
wire		and_181a61d0_u0;
wire		not_141a4211_u0;
wire	[31:0]	mux_19c9b686_u0;
wire		not_494acd65_u0;
reg		done_qual_u135=1'h0;
reg		done_qual_u136_u0=1'h0;
wire		not_256d40f9_u0;
wire		and_5fd20aa7_u0;
reg		done_qual_u137_u0=1'h0;
wire		or_3723931b_u0;
wire	[15:0]	mux_1d7c9d66_u0;
wire		or_26f203ac_u0;
assign and_58fc57bc_u0=or_66105f34_u0&bus_12a00bf7_;
assign or_61208902_u0=bus_4e950722_|done_qual_u136_u0;
assign or_6978c77b_u0=bus_2e13b093_|done_qual_u135;
assign or_66105f34_u0=bus_48029f45_|done_qual_u137_u0;
assign and_181a61d0_u0=or_6978c77b_u0&bus_12a00bf7_;
assign not_141a4211_u0=~bus_12a00bf7_;
assign mux_19c9b686_u0=({32{bus_4e950722_}}&bus_7ccb383c_)|({32{bus_2e13b093_}}&bus_2c80aee2_)|({32{bus_48029f45_}}&bus_0b8f5236_);
assign not_494acd65_u0=~bus_12a00bf7_;
always @(posedge bus_7903d426_)
begin
if (bus_762e0ccd_)
done_qual_u135<=1'h0;
else done_qual_u135<=bus_2e13b093_;
end
assign bus_141e2cb9_=mux_1d7c9d66_u0;
assign bus_62beb692_=mux_19c9b686_u0;
assign bus_4cfcaed6_=or_26f203ac_u0;
assign bus_461cf331_=or_3723931b_u0;
assign bus_5740abcd_=3'h1;
assign bus_402c7489_=and_5fd20aa7_u0;
assign bus_2f4398a5_=and_181a61d0_u0;
assign bus_7b37a050_=bus_0d18c1eb_;
assign bus_43715c56_=and_58fc57bc_u0;
always @(posedge bus_7903d426_)
begin
if (bus_762e0ccd_)
done_qual_u136_u0<=1'h0;
else done_qual_u136_u0<=bus_4e950722_;
end
assign not_256d40f9_u0=~bus_12a00bf7_;
assign and_5fd20aa7_u0=or_61208902_u0&bus_12a00bf7_;
always @(posedge bus_7903d426_)
begin
if (bus_762e0ccd_)
done_qual_u137_u0<=1'h0;
else done_qual_u137_u0<=bus_48029f45_;
end
assign or_3723931b_u0=bus_4e950722_|bus_2e13b093_|bus_48029f45_;
assign mux_1d7c9d66_u0=(bus_4e950722_)?bus_0f7eec10_:bus_75309ed5_;
assign or_26f203ac_u0=bus_4e950722_|bus_2e13b093_;
endmodule



module resized_HH3_xy_endianswapper_3e58fd2a_(endianswapper_3e58fd2a_in, endianswapper_3e58fd2a_out);
input	[31:0]	endianswapper_3e58fd2a_in;
output	[31:0]	endianswapper_3e58fd2a_out;
assign endianswapper_3e58fd2a_out=endianswapper_3e58fd2a_in;
endmodule



module resized_HH3_xy_endianswapper_06a6ceab_(endianswapper_06a6ceab_in, endianswapper_06a6ceab_out);
input	[31:0]	endianswapper_06a6ceab_in;
output	[31:0]	endianswapper_06a6ceab_out;
assign endianswapper_06a6ceab_out=endianswapper_06a6ceab_in;
endmodule



module resized_HH3_xy_stateVar_Out1TokenIndex(bus_1a06ee5a_, bus_21fbc7d7_, bus_11445d5e_, bus_43a7b829_, bus_54879690_);
input		bus_1a06ee5a_;
input		bus_21fbc7d7_;
input		bus_11445d5e_;
input	[31:0]	bus_43a7b829_;
output	[31:0]	bus_54879690_;
wire	[31:0]	endianswapper_3e58fd2a_out;
wire	[31:0]	endianswapper_06a6ceab_out;
reg	[31:0]	stateVar_Out1TokenIndex_u2=32'h0;
resized_HH3_xy_endianswapper_3e58fd2a_ resized_HH3_xy_endianswapper_3e58fd2a__1(.endianswapper_3e58fd2a_in(bus_43a7b829_), 
  .endianswapper_3e58fd2a_out(endianswapper_3e58fd2a_out));
resized_HH3_xy_endianswapper_06a6ceab_ resized_HH3_xy_endianswapper_06a6ceab__1(.endianswapper_06a6ceab_in(stateVar_Out1TokenIndex_u2), 
  .endianswapper_06a6ceab_out(endianswapper_06a6ceab_out));
always @(posedge bus_1a06ee5a_ or posedge bus_21fbc7d7_)
begin
if (bus_21fbc7d7_)
stateVar_Out1TokenIndex_u2<=32'h0;
else if (bus_11445d5e_)
stateVar_Out1TokenIndex_u2<=endianswapper_3e58fd2a_out;
end
assign bus_54879690_=endianswapper_06a6ceab_out;
endmodule



module resized_HH3_xy_simplememoryreferee_233a65d9_(bus_0e63ff2e_, bus_2cbe6427_, bus_0b7a09f9_, bus_3f845529_, bus_51dc5427_, bus_31d29381_, bus_1539b851_, bus_5cf79b2a_, bus_6417eca8_, bus_351c3c2f_, bus_3d2a2664_, bus_27d1116c_, bus_28bc5e54_, bus_1a7956cb_, bus_534cc528_, bus_55d21a89_, bus_4775846d_, bus_0f2a4aab_, bus_7ca17cbb_);
input		bus_0e63ff2e_;
input		bus_2cbe6427_;
input		bus_0b7a09f9_;
input	[15:0]	bus_3f845529_;
input		bus_51dc5427_;
input	[15:0]	bus_31d29381_;
input	[31:0]	bus_1539b851_;
input	[2:0]	bus_5cf79b2a_;
input		bus_6417eca8_;
input	[31:0]	bus_351c3c2f_;
input	[2:0]	bus_3d2a2664_;
output	[15:0]	bus_27d1116c_;
output	[31:0]	bus_28bc5e54_;
output		bus_1a7956cb_;
output		bus_534cc528_;
output	[2:0]	bus_55d21a89_;
output		bus_4775846d_;
output	[15:0]	bus_0f2a4aab_;
output		bus_7ca17cbb_;
wire		not_15983f39_u0;
wire		and_0cb68955_u0;
reg		done_qual_u138_u0=1'h0;
wire	[15:0]	mux_3215a79f_u0;
wire		or_397c15b6_u0;
reg		done_qual_u139_u0=1'h0;
wire		not_6049c599_u0;
wire	[31:0]	mux_7367fdd4_u0;
wire		or_135d7e4e_u0;
wire		or_25c75592_u0;
wire		and_042ac05d_u0;
assign not_15983f39_u0=~bus_0b7a09f9_;
assign and_0cb68955_u0=or_397c15b6_u0&bus_0b7a09f9_;
always @(posedge bus_0e63ff2e_)
begin
if (bus_2cbe6427_)
done_qual_u138_u0<=1'h0;
else done_qual_u138_u0<=bus_51dc5427_;
end
assign mux_3215a79f_u0=({16{bus_51dc5427_}}&bus_31d29381_);
assign or_397c15b6_u0=bus_51dc5427_|done_qual_u138_u0;
always @(posedge bus_0e63ff2e_)
begin
if (bus_2cbe6427_)
done_qual_u139_u0<=1'h0;
else done_qual_u139_u0<=bus_6417eca8_;
end
assign not_6049c599_u0=~bus_0b7a09f9_;
assign mux_7367fdd4_u0=(bus_51dc5427_)?bus_1539b851_:bus_351c3c2f_;
assign or_135d7e4e_u0=bus_51dc5427_|bus_6417eca8_;
assign or_25c75592_u0=bus_6417eca8_|done_qual_u139_u0;
assign and_042ac05d_u0=or_25c75592_u0&bus_0b7a09f9_;
assign bus_27d1116c_=mux_3215a79f_u0;
assign bus_28bc5e54_=mux_7367fdd4_u0;
assign bus_1a7956cb_=bus_51dc5427_;
assign bus_534cc528_=or_135d7e4e_u0;
assign bus_55d21a89_=3'h1;
assign bus_4775846d_=and_0cb68955_u0;
assign bus_0f2a4aab_=bus_3f845529_;
assign bus_7ca17cbb_=and_042ac05d_u0;
endmodule



module resized_HH3_xy_stateVar_Out1PortEnable(bus_4966e2b3_, bus_160bb6e7_, bus_4ad9d6ae_, bus_7fa3f2df_, bus_75e7dd97_);
input		bus_4966e2b3_;
input		bus_160bb6e7_;
input		bus_4ad9d6ae_;
input		bus_7fa3f2df_;
output		bus_75e7dd97_;
reg		stateVar_Out1PortEnable_u2=1'h0;
assign bus_75e7dd97_=stateVar_Out1PortEnable_u2;
always @(posedge bus_4966e2b3_ or posedge bus_160bb6e7_)
begin
if (bus_160bb6e7_)
stateVar_Out1PortEnable_u2<=1'h0;
else if (bus_4ad9d6ae_)
stateVar_Out1PortEnable_u2<=bus_7fa3f2df_;
end
endmodule



module resized_HH3_xy_repeatRowExpanded(CLK, RESET, GO, port_1a399e92_, port_5bdc04de_, port_095c79c5_, port_5a868a9f_, RESULT, RESULT_u1596, RESULT_u1597, RESULT_u1598, RESULT_u1599, RESULT_u1600, RESULT_u1601, RESULT_u1602, RESULT_u1603, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_1a399e92_;
input		port_5bdc04de_;
input	[15:0]	port_095c79c5_;
input		port_5a868a9f_;
output		RESULT;
output	[15:0]	RESULT_u1596;
output		RESULT_u1597;
output	[31:0]	RESULT_u1598;
output	[2:0]	RESULT_u1599;
output		RESULT_u1600;
output	[31:0]	RESULT_u1601;
output	[15:0]	RESULT_u1602;
output	[2:0]	RESULT_u1603;
output		DONE;
wire	[15:0]	add;
wire		and_u2672_u0;
wire		and_u2673_u0;
wire		lessThan;
wire signed	[31:0]	lessThan_b_signed;
wire signed	[31:0]	lessThan_a_signed;
wire		and_u2674_u0;
wire		not_u465_u0;
wire		and_u2675_u0;
reg		and_delayed_u173=1'h0;
wire	[31:0]	add_u269;
wire		and_u2676_u0;
wire	[31:0]	add_u270;
reg		reg_3213c06b_u0=1'h0;
wire		and_u2677_u0;
wire		or_u791_u0;
wire	[31:0]	add_u271;
reg	[31:0]	syncEnable_u433=32'h0;
wire		or_u792_u0;
wire	[31:0]	mux_u269;
reg		reg_39097570_u0=1'h0;
assign add=port_1a399e92_+16'h1;
assign and_u2672_u0=and_u2675_u0&or_u792_u0;
assign and_u2673_u0=and_u2674_u0&or_u792_u0;
assign lessThan_a_signed=mux_u269;
assign lessThan_b_signed=32'h200;
assign lessThan=lessThan_a_signed<lessThan_b_signed;
assign and_u2674_u0=or_u792_u0&not_u465_u0;
assign not_u465_u0=~lessThan;
assign and_u2675_u0=or_u792_u0&lessThan;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u173<=1'h0;
else and_delayed_u173<=and_u2672_u0;
end
assign add_u269=mux_u269+32'h0;
assign and_u2676_u0=and_u2672_u0&port_5bdc04de_;
assign add_u270=mux_u269+32'h0;
always @(posedge CLK or posedge and_u2672_u0 or posedge or_u791_u0)
begin
if (or_u791_u0)
reg_3213c06b_u0<=1'h0;
else if (and_u2672_u0)
reg_3213c06b_u0<=1'h1;
else reg_3213c06b_u0<=reg_3213c06b_u0;
end
assign and_u2677_u0=reg_3213c06b_u0&port_5a868a9f_;
assign or_u791_u0=and_u2677_u0|RESET;
assign add_u271=mux_u269+32'h1;
always @(posedge CLK)
begin
if (and_u2672_u0)
syncEnable_u433<=add_u271;
end
assign or_u792_u0=reg_39097570_u0|and_delayed_u173;
assign mux_u269=(reg_39097570_u0)?32'h0:syncEnable_u433;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_39097570_u0<=1'h0;
else reg_39097570_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u1596=add;
assign RESULT_u1597=and_u2672_u0;
assign RESULT_u1598=add_u269;
assign RESULT_u1599=3'h1;
assign RESULT_u1600=and_u2672_u0;
assign RESULT_u1601=add_u270;
assign RESULT_u1602=port_095c79c5_;
assign RESULT_u1603=3'h1;
assign DONE=and_u2673_u0;
endmodule



module resized_HH3_xy_endianswapper_449152af_(endianswapper_449152af_in, endianswapper_449152af_out);
input	[15:0]	endianswapper_449152af_in;
output	[15:0]	endianswapper_449152af_out;
assign endianswapper_449152af_out=endianswapper_449152af_in;
endmodule



module resized_HH3_xy_endianswapper_5e2d3903_(endianswapper_5e2d3903_in, endianswapper_5e2d3903_out);
input	[15:0]	endianswapper_5e2d3903_in;
output	[15:0]	endianswapper_5e2d3903_out;
assign endianswapper_5e2d3903_out=endianswapper_5e2d3903_in;
endmodule



module resized_HH3_xy_stateVar_x(bus_1f8eca8a_, bus_57b1029e_, bus_0ffcb094_, bus_3935aade_, bus_1fbb8f18_, bus_121158f5_, bus_429824b9_);
input		bus_1f8eca8a_;
input		bus_57b1029e_;
input		bus_0ffcb094_;
input	[15:0]	bus_3935aade_;
input		bus_1fbb8f18_;
input	[15:0]	bus_121158f5_;
output	[15:0]	bus_429824b9_;
wire	[15:0]	mux_0c7481c0_u0;
wire		or_75517448_u0;
reg	[15:0]	stateVar_x_u2=16'h0;
wire	[15:0]	endianswapper_449152af_out;
wire	[15:0]	endianswapper_5e2d3903_out;
assign mux_0c7481c0_u0=(bus_0ffcb094_)?bus_3935aade_:16'h0;
assign or_75517448_u0=bus_0ffcb094_|bus_1fbb8f18_;
always @(posedge bus_1f8eca8a_ or posedge bus_57b1029e_)
begin
if (bus_57b1029e_)
stateVar_x_u2<=16'h0;
else if (or_75517448_u0)
stateVar_x_u2<=endianswapper_449152af_out;
end
assign bus_429824b9_=endianswapper_5e2d3903_out;
resized_HH3_xy_endianswapper_449152af_ resized_HH3_xy_endianswapper_449152af__1(.endianswapper_449152af_in(mux_0c7481c0_u0), 
  .endianswapper_449152af_out(endianswapper_449152af_out));
resized_HH3_xy_endianswapper_5e2d3903_ resized_HH3_xy_endianswapper_5e2d3903__1(.endianswapper_5e2d3903_in(stateVar_x_u2), 
  .endianswapper_5e2d3903_out(endianswapper_5e2d3903_out));
endmodule



module resized_HH3_xy_endianswapper_65a216b4_(endianswapper_65a216b4_in, endianswapper_65a216b4_out);
input		endianswapper_65a216b4_in;
output		endianswapper_65a216b4_out;
assign endianswapper_65a216b4_out=endianswapper_65a216b4_in;
endmodule



module resized_HH3_xy_endianswapper_30f2b1f4_(endianswapper_30f2b1f4_in, endianswapper_30f2b1f4_out);
input		endianswapper_30f2b1f4_in;
output		endianswapper_30f2b1f4_out;
assign endianswapper_30f2b1f4_out=endianswapper_30f2b1f4_in;
endmodule



module resized_HH3_xy_stateVar_fsmState_resized_HH3_xy(bus_49fba71e_, bus_1273375e_, bus_0954f839_, bus_16417063_, bus_5fbc036a_);
input		bus_49fba71e_;
input		bus_1273375e_;
input		bus_0954f839_;
input		bus_16417063_;
output		bus_5fbc036a_;
reg		stateVar_fsmState_resized_HH3_xy_u0=1'h0;
wire		endianswapper_65a216b4_out;
wire		endianswapper_30f2b1f4_out;
always @(posedge bus_49fba71e_ or posedge bus_1273375e_)
begin
if (bus_1273375e_)
stateVar_fsmState_resized_HH3_xy_u0<=1'h0;
else if (bus_0954f839_)
stateVar_fsmState_resized_HH3_xy_u0<=endianswapper_65a216b4_out;
end
resized_HH3_xy_endianswapper_65a216b4_ resized_HH3_xy_endianswapper_65a216b4__1(.endianswapper_65a216b4_in(bus_16417063_), 
  .endianswapper_65a216b4_out(endianswapper_65a216b4_out));
resized_HH3_xy_endianswapper_30f2b1f4_ resized_HH3_xy_endianswapper_30f2b1f4__1(.endianswapper_30f2b1f4_in(stateVar_fsmState_resized_HH3_xy_u0), 
  .endianswapper_30f2b1f4_out(endianswapper_30f2b1f4_out));
assign bus_5fbc036a_=endianswapper_30f2b1f4_out;
endmodule



module resized_HH3_xy_endianswapper_28a9985a_(endianswapper_28a9985a_in, endianswapper_28a9985a_out);
input	[15:0]	endianswapper_28a9985a_in;
output	[15:0]	endianswapper_28a9985a_out;
assign endianswapper_28a9985a_out=endianswapper_28a9985a_in;
endmodule



module resized_HH3_xy_endianswapper_26afe045_(endianswapper_26afe045_in, endianswapper_26afe045_out);
input	[15:0]	endianswapper_26afe045_in;
output	[15:0]	endianswapper_26afe045_out;
assign endianswapper_26afe045_out=endianswapper_26afe045_in;
endmodule



module resized_HH3_xy_stateVar_rowRepeated(bus_003a3253_, bus_7eeb9fab_, bus_0e31d817_, bus_7d7c11ad_, bus_67f23a28_, bus_63962b7e_, bus_1b8c04d2_);
input		bus_003a3253_;
input		bus_7eeb9fab_;
input		bus_0e31d817_;
input	[15:0]	bus_7d7c11ad_;
input		bus_67f23a28_;
input	[15:0]	bus_63962b7e_;
output	[15:0]	bus_1b8c04d2_;
wire	[15:0]	mux_608cdfec_u0;
wire	[15:0]	endianswapper_28a9985a_out;
wire		or_5a6ea134_u0;
wire	[15:0]	endianswapper_26afe045_out;
reg	[15:0]	stateVar_rowRepeated_u2=16'h1;
assign mux_608cdfec_u0=(bus_0e31d817_)?bus_7d7c11ad_:16'h1;
resized_HH3_xy_endianswapper_28a9985a_ resized_HH3_xy_endianswapper_28a9985a__1(.endianswapper_28a9985a_in(mux_608cdfec_u0), 
  .endianswapper_28a9985a_out(endianswapper_28a9985a_out));
assign bus_1b8c04d2_=endianswapper_26afe045_out;
assign or_5a6ea134_u0=bus_0e31d817_|bus_67f23a28_;
resized_HH3_xy_endianswapper_26afe045_ resized_HH3_xy_endianswapper_26afe045__1(.endianswapper_26afe045_in(stateVar_rowRepeated_u2), 
  .endianswapper_26afe045_out(endianswapper_26afe045_out));
always @(posedge bus_003a3253_ or posedge bus_7eeb9fab_)
begin
if (bus_7eeb9fab_)
stateVar_rowRepeated_u2<=16'h1;
else if (or_5a6ea134_u0)
stateVar_rowRepeated_u2<=endianswapper_28a9985a_out;
end
endmodule



module resized_HH3_xy_scheduler(CLK, RESET, GO, port_69930ca0_, port_7545a1a4_, port_1121f1ff_, port_70929f20_, port_05f8f754_, port_697394d7_, port_2ef7caed_, port_1f63f705_, port_0a0e1767_, port_5286b1a6_, port_64176099_, port_21602b46_, port_3915346e_, port_3a6df956_, RESULT, RESULT_u1604, RESULT_u1605, RESULT_u1606, RESULT_u1607, RESULT_u1608, RESULT_u1609, RESULT_u1610, RESULT_u1611, RESULT_u1612, RESULT_u1613, RESULT_u1614, RESULT_u1615, RESULT_u1616, RESULT_u1617, RESULT_u1618, RESULT_u1619, RESULT_u1620, RESULT_u1621, DONE);
input		CLK;
input		RESET;
input		GO;
input	[31:0]	port_69930ca0_;
input		port_7545a1a4_;
input	[31:0]	port_1121f1ff_;
input	[31:0]	port_70929f20_;
input		port_05f8f754_;
input	[15:0]	port_697394d7_;
input	[15:0]	port_2ef7caed_;
input		port_1f63f705_;
input	[15:0]	port_0a0e1767_;
input		port_5286b1a6_;
input		port_64176099_;
input		port_21602b46_;
input		port_3915346e_;
input		port_3a6df956_;
output		RESULT;
output	[31:0]	RESULT_u1604;
output		RESULT_u1605;
output		RESULT_u1606;
output		RESULT_u1607;
output	[31:0]	RESULT_u1608;
output		RESULT_u1609;
output	[31:0]	RESULT_u1610;
output		RESULT_u1611;
output		RESULT_u1612;
output		RESULT_u1613;
output	[31:0]	RESULT_u1614;
output	[2:0]	RESULT_u1615;
output		RESULT_u1616;
output	[15:0]	RESULT_u1617;
output		RESULT_u1618;
output		RESULT_u1619;
output	[15:0]	RESULT_u1620;
output		RESULT_u1621;
output		DONE;
wire	[15:0]	lessThan_b_unsigned;
wire	[15:0]	lessThan_a_unsigned;
wire		lessThan;
wire		equals;
wire	[15:0]	equals_a_unsigned;
wire	[15:0]	equals_b_unsigned;
wire	[15:0]	lessThan_u62_a_unsigned;
wire		lessThan_u62;
wire	[15:0]	lessThan_u62_b_unsigned;
wire		andOp;
wire	[15:0]	equals_u140_b_unsigned;
wire		equals_u140;
wire	[15:0]	equals_u140_a_unsigned;
wire signed	[31:0]	equals_u141_b_signed;
wire signed	[31:0]	equals_u141_a_signed;
wire		equals_u141;
wire		and_u2678_u0;
wire		not_u466_u0;
wire		and_u2679_u0;
wire		andOp_u153;
wire		not_u467_u0;
wire		and_u2680_u0;
wire		and_u2681_u0;
wire		simplePinWrite;
wire		and_u2682_u0;
wire		not_u468_u0;
wire		and_u2683_u0;
wire		simplePinWrite_u416;
wire		not_u469_u0;
wire		and_u2684_u0;
wire		and_u2685_u0;
wire		simplePinWrite_u417;
wire		and_u2686_u0;
reg		reg_3851f050_u0=1'h0;
reg		reg_607d9479_u0=1'h0;
reg		reg_2bfc93f9_u0=1'h0;
reg		reg_23c003c5_u0=1'h0;
reg		reg_38ae08a8_u0=1'h0;
reg		reg_74ed74eb_u0=1'h0;
reg		reg_710aad0d_u0=1'h0;
reg		reg_4cf0ecf8_u0=1'h0;
reg		reg_4cf0ecf8_result_delayed_u0=1'h0;
reg		reg_31f2b9fa_u0=1'h0;
reg		reg_7572dd7f_u0=1'h0;
reg		reg_62f7e6e1_u0=1'h0;
reg		reg_35cd15db_u0=1'h0;
reg		reg_3e561e48_u0=1'h0;
reg		reg_1d95898b_u0=1'h0;
reg		reg_2177b168_u0=1'h0;
reg		reg_3bdd9bc2_u0=1'h0;
reg		reg_459701b4_u0=1'h0;
reg		reg_2d137930_u0=1'h0;
reg		reg_38ae08a8_result_delayed_u0=1'h0;
reg		reg_1d5b7d72_u0=1'h0;
reg		reg_2e8ff2a2_u0=1'h0;
reg		reg_738977bb_u0=1'h0;
reg		reg_47f45fc0_u0=1'h0;
reg		reg_65138d26_u0=1'h0;
reg		reg_12415e78_u0=1'h0;
reg		reg_6a7e8a40_u0=1'h0;
reg		reg_4d591d1c_u0=1'h0;
reg		reg_686a8c2c_u0=1'h0;
reg		reg_6ee35aab_u0=1'h0;
reg		reg_4e9416d8_u0=1'h0;
reg		reg_6c3dc470_u0=1'h0;
reg		reg_4ba6c3eb_u0=1'h0;
reg		reg_4497f4d9_u0=1'h0;
reg		reg_345a7803_u0=1'h0;
reg		reg_1df705ad_u0=1'h0;
reg		reg_5feeefb2_u0=1'h0;
reg		reg_215ed100_u0=1'h0;
reg		reg_4f70c32f_u0=1'h0;
reg		reg_2cc01ca0_u0=1'h0;
reg		reg_5bba6fd9_u0=1'h0;
reg		reg_4e37ba53_u0=1'h0;
reg		reg_01431d27_u0=1'h0;
reg		reg_0e25ee41_u0=1'h0;
reg		reg_051b0973_u0=1'h0;
reg		reg_20d8e0b0_u0=1'h0;
reg		reg_07aa93c1_u0=1'h0;
reg		reg_77c337a8_u0=1'h0;
reg		reg_14095c65_u0=1'h0;
reg		reg_5421084c_u0=1'h0;
reg		reg_33d17fbe_u0=1'h0;
reg		reg_398565f1_u0=1'h0;
reg		reg_2cbb2cce_u0=1'h0;
reg		reg_44757003_u0=1'h0;
reg		reg_098c01f7_u0=1'h0;
reg		reg_7c584cdd_u0=1'h0;
reg		reg_2fda3f5d_u0=1'h0;
reg		reg_46180292_u0=1'h0;
reg		reg_3e132299_u0=1'h0;
reg		reg_6b869f0a_u0=1'h0;
reg		reg_4f7f23f2_u0=1'h0;
reg		reg_133b2fb4_u0=1'h0;
reg		reg_64362ca6_u0=1'h0;
reg		reg_4ecc7e59_u0=1'h0;
reg		reg_3f4f33d9_u0=1'h0;
reg		reg_7399b70f_u0=1'h0;
reg		reg_09c14556_u0=1'h0;
reg		reg_46180292_result_delayed_u0=1'h0;
reg		reg_4e37ba53_result_delayed_u0=1'h0;
reg		reg_46e39e7c_u0=1'h0;
reg		reg_5aa3a23c_u0=1'h0;
reg		reg_6a5362cc_u0=1'h0;
reg		reg_6bfdef5c_u0=1'h0;
reg		reg_4f435be2_u0=1'h0;
reg		reg_686a8c2c_result_delayed_u0=1'h0;
reg		reg_7136b992_u0=1'h0;
reg		reg_30e39c45_u0=1'h0;
reg		reg_2e5316fb_u0=1'h0;
reg		reg_7f08dfa4_u0=1'h0;
reg		reg_0bddd372_u0=1'h0;
reg		reg_35cd15db_result_delayed_u0=1'h0;
reg		reg_39cf897d_u0=1'h0;
reg		reg_42ddc26b_u0=1'h0;
reg		reg_2cf5744d_u0=1'h0;
reg		reg_03c03f7a_u0=1'h0;
reg		reg_1941b9ff_u0=1'h0;
reg		reg_3ddee161_u0=1'h0;
reg		reg_215ed100_result_delayed_u0=1'h0;
reg		reg_3ddee161_result_delayed_u0=1'h0;
wire		or_u793_u0;
reg		reg_357fadb7_u0=1'h0;
reg		reg_02899a41_u0=1'h0;
reg		reg_2cf5703d_u0=1'h0;
reg		reg_5e91ea5a_u0=1'h0;
reg		reg_133b2fb4_result_delayed_u0=1'h0;
reg		reg_3582bd53_u0=1'h0;
reg		reg_33c9371a_u0=1'h0;
reg		reg_7fea3339_u0=1'h0;
reg		reg_328a525c_u0=1'h0;
reg		reg_38c2bc14_u0=1'h0;
reg		reg_0a55fe82_u0=1'h0;
reg		reg_357fadb7_result_delayed_u0=1'h0;
reg		reg_50915049_u0=1'h0;
reg		reg_742b90f1_u0=1'h0;
reg		reg_56c7f61c_u0=1'h0;
reg		reg_377e6fa5_u0=1'h0;
reg		reg_50915049_result_delayed_u0=1'h0;
reg		reg_2cf5703d_result_delayed_u0=1'h0;
reg		reg_42f8ea27_u0=1'h0;
reg		reg_7fea3339_result_delayed_u0=1'h0;
reg		reg_0a125ef3_u0=1'h0;
reg		reg_3ddee161_result_delayed_result_delayed_u0=1'h0;
reg		reg_4f70c32f_result_delayed_u0=1'h0;
reg		reg_67074bef_u0=1'h0;
reg		reg_53cd0b25_u0=1'h0;
reg		reg_4ecc7e59_result_delayed_u0=1'h0;
reg		reg_50915049_result_delayed_result_delayed_u0=1'h0;
reg		reg_47f45fc0_result_delayed_u0=1'h0;
reg		reg_40f72c06_u0=1'h0;
reg		reg_7bbff74c_u0=1'h0;
reg		reg_3dda652e_u0=1'h0;
reg		reg_3fc46730_u0=1'h0;
reg		reg_7f74a383_u0=1'h0;
reg		reg_42ddc26b_result_delayed_u0=1'h0;
reg		reg_4f6a4392_u0=1'h0;
reg		reg_331527ef_u0=1'h0;
reg		reg_1e29aad3_u0=1'h0;
reg		reg_3fd1972f_u0=1'h0;
reg		reg_0ea303a6_u0=1'h0;
wire		and_u2687_u0;
reg		reg_4cade9aa_u0=1'h0;
reg		reg_6052ed5a_u0=1'h0;
reg		reg_5421084c_result_delayed_u0=1'h0;
reg		reg_20d8e0b0_result_delayed_u0=1'h0;
reg		reg_2892d198_u0=1'h0;
reg		reg_23e976e3_u0=1'h0;
reg		reg_07fe52f5_u0=1'h0;
reg		reg_7f74a383_result_delayed_u0=1'h0;
reg		reg_03bbbeb5_u0=1'h0;
reg		reg_00a555b0_u0=1'h0;
reg		reg_16d553cc_u0=1'h0;
reg		reg_45a48cbd_u0=1'h0;
reg		reg_2cf5744d_result_delayed_u0=1'h0;
reg		reg_459701b4_result_delayed_u0=1'h0;
reg		reg_3fd572c8_u0=1'h0;
reg		reg_575abe47_u0=1'h0;
reg		reg_353a7c24_u0=1'h0;
reg		reg_58641d44_u0=1'h0;
reg		reg_6a5362cc_result_delayed_u0=1'h0;
reg		reg_25d144f5_u0=1'h0;
reg		reg_6cdb19fe_u0=1'h0;
reg		reg_6fa4028c_u0=1'h0;
reg		reg_41e078cd_u0=1'h0;
reg		reg_1fd68ee4_u0=1'h0;
reg		reg_7e0acb38_u0=1'h0;
reg		reg_72251f10_u0=1'h0;
reg		reg_2cf5703d_result_delayed_result_delayed_u0=1'h0;
reg		reg_7c7f2949_u0=1'h0;
reg		reg_2cc3d1f5_u0=1'h0;
reg		reg_12fa7fcd_u0=1'h0;
reg		reg_2177b168_result_delayed_u0=1'h0;
reg		reg_2abca780_u0=1'h0;
reg		reg_71dddce1_u0=1'h0;
reg		reg_4d587466_u0=1'h0;
reg		reg_72076745_u0=1'h0;
reg		reg_6ff6deb2_u0=1'h0;
reg		reg_3d9590d0_u0=1'h0;
reg		reg_01f5f8bd_u0=1'h0;
reg		reg_1a8e23c7_u0=1'h0;
reg		reg_7ab59fff_u0=1'h0;
reg		reg_4e37ba53_result_delayed_result_delayed_u0=1'h0;
reg		reg_7bbff74c_result_delayed_u0=1'h0;
reg		reg_77c337a8_result_delayed_u0=1'h0;
reg		reg_2892d198_result_delayed_u0=1'h0;
reg		reg_6b869f0a_result_delayed_u0=1'h0;
reg		reg_2db318e2_u0=1'h0;
reg		reg_57c45696_u0=1'h0;
reg		reg_658e74db_u0=1'h0;
reg		reg_38c2bc14_result_delayed_u0=1'h0;
reg		reg_4b8c12d0_u0=1'h0;
reg		reg_01347069_u0=1'h0;
reg		reg_4e37ba53_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_328a525c_result_delayed_u0=1'h0;
reg		reg_2cc3d1f5_result_delayed_u0=1'h0;
reg		reg_1c090d6c_u0=1'h0;
reg		reg_33c9371a_result_delayed_u0=1'h0;
reg		reg_3851f050_result_delayed_u0=1'h0;
reg		reg_2e8ff2a2_result_delayed_u0=1'h0;
reg		reg_0414817f_u0=1'h0;
reg		reg_185bb135_u0=1'h0;
reg		reg_1b3d5a52_u0=1'h0;
reg		reg_2c350944_u0=1'h0;
reg		reg_2af4ab86_u0=1'h0;
reg		reg_3113d461_u0=1'h0;
reg		reg_295e5824_u0=1'h0;
reg		reg_46180292_result_delayed_result_delayed_u0=1'h0;
reg		reg_38ae08a8_result_delayed_result_delayed_u0=1'h0;
reg		reg_5e62c71d_u0=1'h0;
reg		reg_44757003_result_delayed_u0=1'h0;
reg		reg_7136b992_result_delayed_u0=1'h0;
reg		reg_53b43e36_u0=1'h0;
reg		reg_377e6fa5_result_delayed_u0=1'h0;
reg		reg_7ac1bb42_u0=1'h0;
reg		reg_7fd56e50_u0=1'h0;
reg		reg_119a281f_u0=1'h0;
reg		reg_119a281f_result_delayed_u0=1'h0;
reg		reg_030ef688_u0=1'h0;
reg		reg_42ddc26b_result_delayed_result_delayed_u0=1'h0;
reg		reg_13f4d67d_u0=1'h0;
reg		reg_5fbaaa33_u0=1'h0;
reg		reg_032d42a6_u0=1'h0;
reg		reg_5dc60849_u0=1'h0;
reg		reg_571dd692_u0=1'h0;
reg		reg_4ba6c3eb_result_delayed_u0=1'h0;
reg		reg_382559bf_u0=1'h0;
reg		reg_19da6841_u0=1'h0;
reg		reg_7d04d098_u0=1'h0;
reg		reg_6ee35aab_result_delayed_u0=1'h0;
reg		reg_7d04d098_result_delayed_u0=1'h0;
reg		reg_0ef27753_u0=1'h0;
reg		reg_6ff6deb2_result_delayed_u0=1'h0;
reg		reg_1d5b7d72_result_delayed_u0=1'h0;
reg		reg_2defdc44_u0=1'h0;
reg		reg_5bba6fd9_result_delayed_u0=1'h0;
reg		reg_01f5f8bd_result_delayed_u0=1'h0;
reg		reg_6d8ffc20_u0=1'h0;
reg		reg_6cdb19fe_result_delayed_u0=1'h0;
reg		reg_7f74a383_result_delayed_result_delayed_u0=1'h0;
reg		reg_735e96ed_u0=1'h0;
reg		reg_6bf27e46_u0=1'h0;
reg		reg_5c28119c_u0=1'h0;
reg		reg_07aa93c1_result_delayed_u0=1'h0;
reg		reg_072c9294_u0=1'h0;
reg		reg_5091952b_u0=1'h0;
reg		reg_7ce31523_u0=1'h0;
reg		reg_25d144f5_result_delayed_u0=1'h0;
reg		reg_12415e78_result_delayed_u0=1'h0;
reg		reg_35cd15db_result_delayed_result_delayed_u0=1'h0;
reg		reg_40f72c06_result_delayed_u0=1'h0;
reg		reg_3e561e48_result_delayed_u0=1'h0;
reg		reg_57c45696_result_delayed_u0=1'h0;
reg		reg_6a6f9fa5_u0=1'h0;
reg		reg_7c87d14d_u0=1'h0;
reg		reg_0ef27753_result_delayed_u0=1'h0;
reg		reg_00a555b0_result_delayed_u0=1'h0;
reg		reg_1941b9ff_result_delayed_u0=1'h0;
reg		reg_28b4d165_u0=1'h0;
reg		reg_15ccc01d_u0=1'h0;
reg		reg_2cc3d1f5_result_delayed_result_delayed_u0=1'h0;
reg		reg_09c14556_result_delayed_u0=1'h0;
reg		reg_32854b5c_u0=1'h0;
reg		reg_6134ccef_u0=1'h0;
reg		reg_7572dd7f_result_delayed_u0=1'h0;
reg		reg_30e39c45_result_delayed_u0=1'h0;
reg		reg_6ed66f32_u0=1'h0;
reg		reg_78342dd1_u0=1'h0;
reg		reg_0f9d1678_u0=1'h0;
reg		reg_0414817f_result_delayed_u0=1'h0;
reg		reg_4f852262_u0=1'h0;
reg		reg_023bffd6_u0=1'h0;
reg		reg_596f7c82_u0=1'h0;
reg		reg_6ca72548_u0=1'h0;
reg		reg_1fd68ee4_result_delayed_u0=1'h0;
reg		reg_07fe52f5_result_delayed_u0=1'h0;
reg		reg_16d553cc_result_delayed_u0=1'h0;
reg		reg_1b102eec_u0=1'h0;
reg		reg_63f53a08_u0=1'h0;
reg		reg_38ae08a8_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_4cade9aa_result_delayed_u0=1'h0;
reg		reg_795d0757_u0=1'h0;
reg		reg_44757003_result_delayed_result_delayed_u0=1'h0;
reg		reg_751aa708_u0=1'h0;
reg		reg_1479ea6c_u0=1'h0;
reg		reg_33c9371a_result_delayed_result_delayed_u0=1'h0;
reg		reg_3e2b8c33_u0=1'h0;
reg		reg_2af4ab86_result_delayed_u0=1'h0;
reg		reg_1941b9ff_result_delayed_result_delayed_u0=1'h0;
reg		reg_250a9f11_u0=1'h0;
reg		reg_7b11510d_u0=1'h0;
reg		reg_4497f4d9_result_delayed_u0=1'h0;
reg		reg_39cf897d_result_delayed_u0=1'h0;
reg		reg_0054d249_u0=1'h0;
reg		reg_74ed74eb_result_delayed_u0=1'h0;
reg		reg_2b8f21ae_u0=1'h0;
reg		reg_1f57f175_u0=1'h0;
reg		reg_28b4d165_result_delayed_u0=1'h0;
reg		reg_2e407063_u0=1'h0;
reg		reg_0e5cbc7b_u0=1'h0;
reg		reg_5b704959_u0=1'h0;
reg		reg_4f7f23f2_result_delayed_u0=1'h0;
reg		reg_6ed66f32_result_delayed_u0=1'h0;
reg		reg_357fadb7_result_delayed_result_delayed_u0=1'h0;
reg		reg_03bbbeb5_result_delayed_u0=1'h0;
reg		reg_2be729d4_u0=1'h0;
reg		reg_63f53a08_result_delayed_u0=1'h0;
reg		reg_4e6c385a_u0=1'h0;
reg		reg_0bddd372_result_delayed_u0=1'h0;
reg		reg_2cf5744d_result_delayed_result_delayed_u0=1'h0;
reg		reg_0576bf35_u0=1'h0;
reg		reg_33d17fbe_result_delayed_u0=1'h0;
reg		reg_14095c65_result_delayed_u0=1'h0;
reg		reg_46e39e7c_result_delayed_u0=1'h0;
reg		reg_2cc01ca0_result_delayed_u0=1'h0;
reg		reg_7ac1bb42_result_delayed_u0=1'h0;
reg		reg_4d587466_result_delayed_u0=1'h0;
reg		reg_45a48cbd_result_delayed_u0=1'h0;
reg		reg_2cfcc2a4_u0=1'h0;
reg		reg_43fabda0_u0=1'h0;
reg		reg_79022b5e_u0=1'h0;
reg		reg_3fc46730_result_delayed_u0=1'h0;
reg		reg_35cd15db_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_2a22ac7d_u0=1'h0;
reg		reg_3893a2cc_u0=1'h0;
reg		reg_55043b64_u0=1'h0;
reg		reg_6134ccef_result_delayed_u0=1'h0;
wire		and_u2688_u0;
reg		reg_58980aff_u0=1'h0;
reg		reg_3156ef3e_u0=1'h0;
reg		reg_5feeefb2_result_delayed_u0=1'h0;
reg		reg_14905eff_u0=1'h0;
reg		reg_03bbbeb5_result_delayed_result_delayed_u0=1'h0;
reg		reg_07fe52f5_result_delayed_result_delayed_u0=1'h0;
reg		reg_0576bf35_result_delayed_u0=1'h0;
reg		reg_30e39c45_result_delayed_result_delayed_u0=1'h0;
reg		reg_3843f63d_u0=1'h0;
reg		reg_01f5f8bd_result_delayed_result_delayed_u0=1'h0;
reg		reg_2be729d4_result_delayed_u0=1'h0;
reg		reg_79022b5e_result_delayed_u0=1'h0;
reg		reg_23e976e3_result_delayed_u0=1'h0;
reg		reg_790c1f8e_u0=1'h0;
reg		reg_47f45fc0_result_delayed_result_delayed_u0=1'h0;
reg		reg_217203f5_u0=1'h0;
reg		reg_6aa4982f_u0=1'h0;
reg		reg_16d553cc_result_delayed_result_delayed_u0=1'h0;
reg		reg_795d0757_result_delayed_u0=1'h0;
reg		reg_2cf5744d_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_4f70c32f_result_delayed_result_delayed_u0=1'h0;
reg		reg_2e5316fb_result_delayed_u0=1'h0;
reg		reg_04fc925c_u0=1'h0;
reg		reg_62f7e6e1_result_delayed_u0=1'h0;
reg		reg_710aad0d_result_delayed_u0=1'h0;
reg		reg_32854b5c_result_delayed_u0=1'h0;
reg		reg_1d95898b_result_delayed_u0=1'h0;
reg		reg_25d144f5_result_delayed_result_delayed_u0=1'h0;
reg		reg_686a8c2c_result_delayed_result_delayed_u0=1'h0;
reg		reg_058dcb20_u0=1'h0;
reg		reg_5bba6fd9_result_delayed_result_delayed_u0=1'h0;
reg		reg_43fabda0_result_delayed_u0=1'h0;
reg		reg_4f70c32f_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_5574bbc5_u0=1'h0;
reg		reg_607d9479_result_delayed_u0=1'h0;
reg		reg_3fd1972f_result_delayed_u0=1'h0;
reg		reg_38ae08a8_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_6c3dc470_result_delayed_u0=1'h0;
reg		reg_0b346188_u0=1'h0;
reg		reg_38ae08a8_result_delayed_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_7572dd7f_result_delayed_result_delayed_u0=1'h0;
reg		reg_75d7ab69_u0=1'h0;
reg		reg_1d65b7da_u0=1'h0;
reg		reg_1eed982d_u0=1'h0;
reg		reg_1479ea6c_result_delayed_u0=1'h0;
reg		reg_42f8ea27_result_delayed_u0=1'h0;
reg		reg_4a16e8d3_u0=1'h0;
reg		reg_2cf5744d_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_2be729d4_result_delayed_result_delayed_u0=1'h0;
reg		reg_3893a2cc_result_delayed_u0=1'h0;
reg		reg_5aa3a23c_result_delayed_u0=1'h0;
reg		reg_051b0973_result_delayed_u0=1'h0;
reg		reg_331527ef_result_delayed_u0=1'h0;
reg		reg_01347069_result_delayed_u0=1'h0;
reg		reg_3fd572c8_result_delayed_u0=1'h0;
reg		reg_20d8e0b0_result_delayed_result_delayed_u0=1'h0;
reg		reg_12415e78_result_delayed_result_delayed_u0=1'h0;
reg		reg_6d8ffc20_result_delayed_u0=1'h0;
reg		reg_738977bb_result_delayed_u0=1'h0;
reg		reg_6ff6deb2_result_delayed_result_delayed_u0=1'h0;
reg		reg_658e74db_result_delayed_u0=1'h0;
reg		reg_5d8a9f60_u0=1'h0;
reg		reg_30e39c45_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_023bffd6_result_delayed_u0=1'h0;
reg		reg_4e9416d8_result_delayed_u0=1'h0;
reg		reg_27aff15e_u0=1'h0;
reg		reg_331527ef_result_delayed_result_delayed_u0=1'h0;
reg		reg_30e39c45_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_353a7c24_result_delayed_u0=1'h0;
reg		reg_5d8a9f60_result_delayed_u0=1'h0;
reg		reg_2892d198_result_delayed_result_delayed_u0=1'h0;
reg		reg_2cbb2cce_result_delayed_u0=1'h0;
reg		reg_7136b992_result_delayed_result_delayed_u0=1'h0;
reg		reg_133b2fb4_result_delayed_result_delayed_u0=1'h0;
reg		reg_0a55fe82_result_delayed_u0=1'h0;
reg		reg_2892d198_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_7b11510d_result_delayed_u0=1'h0;
reg		reg_795d0757_result_delayed_result_delayed_u0=1'h0;
reg		reg_0e5cbc7b_result_delayed_u0=1'h0;
reg		reg_5421084c_result_delayed_result_delayed_u0=1'h0;
reg		reg_7c584cdd_result_delayed_u0=1'h0;
reg		reg_571dd692_result_delayed_u0=1'h0;
reg		reg_575abe47_result_delayed_u0=1'h0;
reg		reg_12fa7fcd_result_delayed_u0=1'h0;
reg		reg_331527ef_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_38ae08a8_result_delayed_result_delayed_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_658e74db_result_delayed_result_delayed_u0=1'h0;
reg		reg_6761984a_u0=1'h0;
reg		reg_0963c64e_u0=1'h0;
reg		reg_3f4f33d9_result_delayed_u0=1'h0;
reg		reg_751aa708_result_delayed_u0=1'h0;
reg		reg_4ecc7e59_result_delayed_result_delayed_u0=1'h0;
reg		reg_2a4e2976_u0=1'h0;
reg		reg_0b46a87d_u0=1'h0;
reg		reg_1eed982d_result_delayed_u0=1'h0;
reg		reg_6ed66f32_result_delayed_result_delayed_u0=1'h0;
reg		reg_3113d461_result_delayed_u0=1'h0;
reg		reg_3851f050_result_delayed_result_delayed_u0=1'h0;
reg		reg_67074bef_result_delayed_u0=1'h0;
reg		reg_5b704959_result_delayed_u0=1'h0;
reg		reg_05509604_u0=1'h0;
reg		reg_3582bd53_result_delayed_u0=1'h0;
wire		or_u794_u0;
wire		mux_u270;
reg		reg_46180292_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_2e5316fb_result_delayed_result_delayed_u0=1'h0;
reg		reg_46180292_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_1b102eec_result_delayed_u0=1'h0;
reg		reg_39cf897d_result_delayed_result_delayed_u0=1'h0;
reg		reg_459701b4_result_delayed_result_delayed_u0=1'h0;
reg		reg_6ff6deb2_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_7d04d098_result_delayed_result_delayed_u0=1'h0;
reg		reg_58980aff_result_delayed_u0=1'h0;
reg		reg_7399b70f_result_delayed_u0=1'h0;
reg		reg_4ba6c3eb_result_delayed_result_delayed_u0=1'h0;
reg		reg_3bdd9bc2_result_delayed_u0=1'h0;
reg		reg_2a4e2976_result_delayed_u0=1'h0;
reg		reg_382559bf_result_delayed_u0=1'h0;
reg		reg_7fea3339_result_delayed_result_delayed_u0=1'h0;
reg		reg_32854b5c_result_delayed_result_delayed_u0=1'h0;
reg		reg_75d7ab69_result_delayed_u0=1'h0;
reg		reg_4497f4d9_result_delayed_result_delayed_u0=1'h0;
reg		reg_4f435be2_result_delayed_u0=1'h0;
reg		reg_0f9d1678_result_delayed_u0=1'h0;
reg		reg_7fd56e50_result_delayed_u0=1'h0;
reg		reg_3e132299_result_delayed_u0=1'h0;
reg		reg_2e5316fb_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_098c01f7_result_delayed_u0=1'h0;
reg		reg_032d42a6_result_delayed_u0=1'h0;
reg		reg_65138d26_result_delayed_u0=1'h0;
reg		reg_57c45696_result_delayed_result_delayed_u0=1'h0;
reg		reg_742b90f1_result_delayed_u0=1'h0;
reg		reg_78342dd1_result_delayed_u0=1'h0;
reg		reg_2bfc93f9_result_delayed_u0=1'h0;
reg		reg_6b869f0a_result_delayed_result_delayed_u0=1'h0;
reg		reg_0576bf35_result_delayed_result_delayed_u0=1'h0;
reg		reg_0576bf35_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_7c7f2949_result_delayed_u0=1'h0;
reg		reg_3cf3ff64_u0=1'h0;
reg		reg_185bb135_result_delayed_u0=1'h0;
reg		reg_7b11510d_result_delayed_result_delayed_u0=1'h0;
reg		reg_3bdd9bc2_result_delayed_result_delayed_u0=1'h0;
reg		reg_1d65b7da_result_delayed_u0=1'h0;
reg		reg_398565f1_result_delayed_u0=1'h0;
reg		reg_6ca72548_result_delayed_u0=1'h0;
reg		reg_345a7803_result_delayed_u0=1'h0;
reg		reg_5d8a9f60_result_delayed_result_delayed_u0=1'h0;
reg		reg_571dd692_result_delayed_result_delayed_u0=1'h0;
reg		reg_328a525c_result_delayed_result_delayed_u0=1'h0;
reg		reg_0a125ef3_result_delayed_u0=1'h0;
reg		reg_3cf3ff64_result_delayed_u0=1'h0;
reg		reg_4b4698ef_u0=1'h0;
reg		reg_07aa93c1_result_delayed_result_delayed_u0=1'h0;
reg		reg_0e5cbc7b_result_delayed_result_delayed_u0=1'h0;
reg		reg_14905eff_result_delayed_u0=1'h0;
reg		reg_051b0973_result_delayed_result_delayed_u0=1'h0;
reg		reg_1df705ad_result_delayed_u0=1'h0;
reg		reg_3dda652e_result_delayed_u0=1'h0;
reg		reg_2fda3f5d_result_delayed_u0=1'h0;
reg		reg_1479ea6c_result_delayed_result_delayed_u0=1'h0;
reg		reg_217203f5_result_delayed_u0=1'h0;
reg		reg_1d95898b_result_delayed_result_delayed_u0=1'h0;
reg		reg_2a22ac7d_result_delayed_u0=1'h0;
reg		reg_2f3b2083_u0=1'h0;
reg		reg_31f2b9fa_result_delayed_u0=1'h0;
reg		reg_119a281f_result_delayed_result_delayed_u0=1'h0;
reg		reg_43fabda0_result_delayed_result_delayed_u0=1'h0;
reg		reg_31f2b9fa_result_delayed_result_delayed_u0=1'h0;
reg		reg_795d0757_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_6134ccef_result_delayed_result_delayed_u0=1'h0;
reg		reg_77c337a8_result_delayed_result_delayed_u0=1'h0;
reg		reg_71dddce1_result_delayed_u0=1'h0;
reg		reg_2f3b2083_result_delayed_u0=1'h0;
reg		reg_7ce31523_result_delayed_u0=1'h0;
reg		reg_459701b4_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_09485a92_u0=1'h0;
reg		reg_3843f63d_result_delayed_u0=1'h0;
reg		reg_0ef27753_result_delayed_result_delayed_u0=1'h0;
reg		reg_23c003c5_result_delayed_u0=1'h0;
reg		reg_4f70c32f_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_2cc01ca0_result_delayed_result_delayed_u0=1'h0;
reg		reg_3582bd53_result_delayed_result_delayed_u0=1'h0;
reg		reg_1a8e23c7_result_delayed_u0=1'h0;
reg		reg_0b346188_result_delayed_u0=1'h0;
reg		reg_11bf5a5d_u0=1'h0;
reg		reg_7b11510d_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_16d553cc_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_4cf0ecf8_result_delayed_result_delayed_u0=1'h0;
reg		reg_46180292_result_delayed_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_1d5b7d72_result_delayed_result_delayed_u0=1'h0;
reg		reg_2892d198_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_33d17fbe_result_delayed_result_delayed_u0=1'h0;
reg		reg_7bbff74c_result_delayed_result_delayed_u0=1'h0;
reg		reg_4d591d1c_result_delayed_u0=1'h0;
reg		and_delayed_u174=1'h0;
reg		reg_2c350944_result_delayed_u0=1'h0;
reg		reg_6ff6deb2_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_2d137930_result_delayed_u0=1'h0;
reg		reg_42f8ea27_result_delayed_result_delayed_u0=1'h0;
reg		reg_0a55fe82_result_delayed_result_delayed_u0=1'h0;
reg		reg_55043b64_result_delayed_u0=1'h0;
reg		reg_50915049_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_7c87d14d_result_delayed_u0=1'h0;
reg		reg_0c581759_u0=1'h0;
reg		reg_3fcc3d8e_u0=1'h0;
wire		or_u795_u0;
wire		or_u796_u0;
wire		or_u797_u0;
wire		or_u798_u0;
reg		reg_102f357e_u0=1'h0;
reg		reg_7b7cf4e5_u0=1'h0;
wire		and_u2689_u0;
reg		reg_0c581759_result_delayed_u0=1'h0;
reg		reg_3fcc3d8e_result_delayed_u0=1'h0;
wire		and_u2690_u0;
reg		reg_102f357e_result_delayed_u0=1'h0;
wire		or_u799_u0;
wire		mux_u271_u0;
reg		reg_0c581759_result_delayed_result_delayed_u0=1'h0;
wire		or_u800_u0;
wire	[31:0]	mux_u272_u0;
reg		reg_102f357e_result_delayed_result_delayed_u0=1'h0;
wire		and_u2691_u0;
reg		reg_6e7913b6_u0=1'h0;
wire		or_u801_u0;
wire		and_u2692_u0;
wire signed	[31:0]	equals_u142_b_signed;
wire signed	[31:0]	equals_u142_a_signed;
wire		equals_u142;
wire		not_u470_u0;
wire		and_u2693_u0;
wire		and_u2694_u0;
wire		and_u2695_u0;
wire		and_u2696_u0;
wire		not_u471_u0;
wire		lessThan_u63;
wire signed	[31:0]	lessThan_u63_b_signed;
wire signed	[31:0]	lessThan_u63_a_signed;
wire		and_u2697_u0;
wire		not_u472_u0;
wire		and_u2698_u0;
wire		not_u473_u0;
wire		and_u2699_u0;
wire		and_u2700_u0;
wire	[31:0]	add;
wire		and_u2701_u0;
wire	[15:0]	simplePinWrite_u418;
wire		simplePinWrite_u419;
wire	[15:0]	simplePinWrite_u420;
wire	[31:0]	add_u272;
reg	[15:0]	syncEnable_u434=16'h0;
reg	[15:0]	syncEnable_u435_u0=16'h0;
wire		and_u2702_u0;
wire		and_u2703_u0;
wire	[15:0]	mux_u273_u0;
reg		and_delayed_u175_u0=1'h0;
reg		and_delayed_u176_u0=1'h0;
reg		reg_0f183598_u0=1'h0;
reg		reg_4418b1bb_u0=1'h0;
wire	[31:0]	mux_u274_u0;
reg	[31:0]	syncEnable_u436_u0=32'h0;
wire		and_u2704_u0;
reg	[15:0]	syncEnable_u437_u0=16'h0;
wire	[15:0]	mux_u275_u0;
wire		and_u2705_u0;
reg		reg_532d6b49_u0=1'h0;
reg		reg_0b4f0828_u0=1'h0;
reg	[31:0]	syncEnable_u438_u0=32'h0;
wire	[15:0]	mux_u276_u0;
reg	[15:0]	syncEnable_u439_u0=16'h0;
wire	[31:0]	mux_u277_u0;
wire		and_u2706_u0;
wire		and_u2707_u0;
wire		and_u2708_u0;
reg		reg_67514dd2_u0=1'h0;
wire	[31:0]	mux_u278_u0;
wire	[15:0]	mux_u279_u0;
reg	[31:0]	syncEnable_u440_u0=32'h0;
wire		and_u2709_u0;
reg	[15:0]	syncEnable_u441_u0=16'h0;
reg		and_delayed_u177_u0=1'h0;
reg		block_GO_delayed_u9=1'h0;
wire		mux_u280_u0;
wire		or_u802_u0;
wire	[31:0]	latch_06dfa717_out;
reg	[31:0]	latch_06dfa717_reg=32'h0;
reg	[15:0]	latch_577ad7b1_reg=16'h0;
wire	[15:0]	latch_577ad7b1_out;
wire	[31:0]	mux_u281_u0;
wire		or_u803_u0;
wire		or_u804_u0;
wire		mux_u282_u0;
wire		or_u805_u0;
wire	[31:0]	mux_u283_u0;
wire		and_u2710_u0;
reg	[31:0]	fbReg_temp_fsmOldState_resized_HH3_xy_5_u0=32'h0;
wire	[15:0]	mux_u284_u0;
reg		syncEnable_u442_u0=1'h0;
reg	[15:0]	fbReg_Out1Portvalue_u2=16'h0;
wire		or_u806_u0;
wire	[31:0]	mux_u285_u0;
reg		loopControl_u6=1'h0;
reg		reg_6f91e613_u0=1'h0;
wire	[31:0]	mux_u286_u0;
wire		or_u807_u0;
wire		or_u808_u0;
wire	[31:0]	mux_u287_u0;
reg		reg_6f91e613_result_delayed_u0=1'h0;
wire		or_u809_u0;
wire		mux_u288_u0;
wire		or_u810_u0;
wire		mux_u289_u0;
wire		or_u811_u0;
assign lessThan_a_unsigned=port_697394d7_;
assign lessThan_b_unsigned=16'h40;
assign lessThan=lessThan_a_unsigned<lessThan_b_unsigned;
assign equals_a_unsigned=port_697394d7_;
assign equals_b_unsigned=16'h40;
assign equals=equals_a_unsigned==equals_b_unsigned;
assign lessThan_u62_a_unsigned=port_2ef7caed_;
assign lessThan_u62_b_unsigned=16'h8;
assign lessThan_u62=lessThan_u62_a_unsigned<lessThan_u62_b_unsigned;
assign andOp=equals&lessThan_u62;
assign equals_u140_a_unsigned=port_2ef7caed_;
assign equals_u140_b_unsigned=16'h8;
assign equals_u140=equals_u140_a_unsigned==equals_u140_b_unsigned;
assign equals_u141_a_signed={31'b0, port_7545a1a4_};
assign equals_u141_b_signed=32'h0;
assign equals_u141=equals_u141_a_signed==equals_u141_b_signed;
assign and_u2678_u0=and_u2710_u0&equals_u141;
assign not_u466_u0=~equals_u141;
assign and_u2679_u0=and_u2710_u0&not_u466_u0;
assign andOp_u153=lessThan&port_21602b46_;
assign not_u467_u0=~andOp_u153;
assign and_u2680_u0=and_u2691_u0&not_u467_u0;
assign and_u2681_u0=and_u2691_u0&andOp_u153;
assign simplePinWrite=and_u2690_u0&{1{and_u2690_u0}};
assign and_u2682_u0=and_u2689_u0&andOp;
assign not_u468_u0=~andOp;
assign and_u2683_u0=and_u2689_u0&not_u468_u0;
assign simplePinWrite_u416=and_u2687_u0&{1{and_u2687_u0}};
assign not_u469_u0=~equals_u140;
assign and_u2684_u0=and_u2688_u0&not_u469_u0;
assign and_u2685_u0=and_u2688_u0&equals_u140;
assign simplePinWrite_u417=and_u2686_u0&{1{and_u2686_u0}};
assign and_u2686_u0=and_u2685_u0&and_u2688_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3851f050_u0<=1'h0;
else reg_3851f050_u0<=reg_6a7e8a40_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_607d9479_u0<=1'h0;
else reg_607d9479_u0<=reg_1fd68ee4_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2bfc93f9_u0<=1'h0;
else reg_2bfc93f9_u0<=reg_6ed66f32_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_23c003c5_u0<=1'h0;
else reg_23c003c5_u0<=reg_04fc925c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_38ae08a8_u0<=1'h0;
else reg_38ae08a8_u0<=reg_78342dd1_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_74ed74eb_u0<=1'h0;
else reg_74ed74eb_u0<=reg_4b4698ef_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_710aad0d_u0<=1'h0;
else reg_710aad0d_u0<=reg_01431d27_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4cf0ecf8_u0<=1'h0;
else reg_4cf0ecf8_u0<=reg_00a555b0_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4cf0ecf8_result_delayed_u0<=1'h0;
else reg_4cf0ecf8_result_delayed_u0<=reg_4cf0ecf8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_31f2b9fa_u0<=1'h0;
else reg_31f2b9fa_u0<=reg_742b90f1_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7572dd7f_u0<=1'h0;
else reg_7572dd7f_u0<=reg_03c03f7a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_62f7e6e1_u0<=1'h0;
else reg_62f7e6e1_u0<=reg_14095c65_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_35cd15db_u0<=1'h0;
else reg_35cd15db_u0<=reg_2cf5703d_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3e561e48_u0<=1'h0;
else reg_3e561e48_u0<=reg_4f6a4392_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1d95898b_u0<=1'h0;
else reg_1d95898b_u0<=reg_1e29aad3_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2177b168_u0<=1'h0;
else reg_2177b168_u0<=reg_030ef688_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3bdd9bc2_u0<=1'h0;
else reg_3bdd9bc2_u0<=reg_7136b992_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_459701b4_u0<=1'h0;
else reg_459701b4_u0<=reg_19da6841_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2d137930_u0<=1'h0;
else reg_2d137930_u0<=reg_058dcb20_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_38ae08a8_result_delayed_u0<=1'h0;
else reg_38ae08a8_result_delayed_u0<=reg_38ae08a8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1d5b7d72_u0<=1'h0;
else reg_1d5b7d72_u0<=reg_0414817f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2e8ff2a2_u0<=1'h0;
else reg_2e8ff2a2_u0<=reg_7f08dfa4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_738977bb_u0<=1'h0;
else reg_738977bb_u0<=reg_50915049_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_47f45fc0_u0<=1'h0;
else reg_47f45fc0_u0<=reg_5574bbc5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_65138d26_u0<=1'h0;
else reg_65138d26_u0<=reg_5e62c71d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_12415e78_u0<=1'h0;
else reg_12415e78_u0<=reg_596f7c82_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6a7e8a40_u0<=1'h0;
else reg_6a7e8a40_u0<=reg_2f3b2083_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4d591d1c_u0<=1'h0;
else reg_4d591d1c_u0<=reg_4f435be2_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_686a8c2c_u0<=1'h0;
else reg_686a8c2c_u0<=reg_1c090d6c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6ee35aab_u0<=1'h0;
else reg_6ee35aab_u0<=reg_5bba6fd9_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4e9416d8_u0<=1'h0;
else reg_4e9416d8_u0<=reg_215ed100_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6c3dc470_u0<=1'h0;
else reg_6c3dc470_u0<=reg_3d9590d0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4ba6c3eb_u0<=1'h0;
else reg_4ba6c3eb_u0<=reg_0e25ee41_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4497f4d9_u0<=1'h0;
else reg_4497f4d9_u0<=reg_3ddee161_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_345a7803_u0<=1'h0;
else reg_345a7803_u0<=reg_2cfcc2a4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1df705ad_u0<=1'h0;
else reg_1df705ad_u0<=reg_4f852262_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5feeefb2_u0<=1'h0;
else reg_5feeefb2_u0<=reg_0576bf35_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_215ed100_u0<=1'h0;
else reg_215ed100_u0<=reg_6a6f9fa5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4f70c32f_u0<=1'h0;
else reg_4f70c32f_u0<=and_u2687_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2cc01ca0_u0<=1'h0;
else reg_2cc01ca0_u0<=reg_3156ef3e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5bba6fd9_u0<=1'h0;
else reg_5bba6fd9_u0<=reg_3f4f33d9_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4e37ba53_u0<=1'h0;
else reg_4e37ba53_u0<=reg_58980aff_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01431d27_u0<=1'h0;
else reg_01431d27_u0<=reg_2af4ab86_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0e25ee41_u0<=1'h0;
else reg_0e25ee41_u0<=reg_32854b5c_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_051b0973_u0<=1'h0;
else reg_051b0973_u0<=reg_4e37ba53_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_20d8e0b0_u0<=1'h0;
else reg_20d8e0b0_u0<=reg_28b4d165_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_07aa93c1_u0<=1'h0;
else reg_07aa93c1_u0<=reg_16d553cc_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_77c337a8_u0<=1'h0;
else reg_77c337a8_u0<=reg_2cc3d1f5_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_14095c65_u0<=1'h0;
else reg_14095c65_u0<=reg_23c003c5_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5421084c_u0<=1'h0;
else reg_5421084c_u0<=reg_6052ed5a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_33d17fbe_u0<=1'h0;
else reg_33d17fbe_u0<=reg_6bfdef5c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_398565f1_u0<=1'h0;
else reg_398565f1_u0<=reg_09c14556_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2cbb2cce_u0<=1'h0;
else reg_2cbb2cce_u0<=reg_098c01f7_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_44757003_u0<=1'h0;
else reg_44757003_u0<=reg_64362ca6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_098c01f7_u0<=1'h0;
else reg_098c01f7_u0<=reg_7e0acb38_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7c584cdd_u0<=1'h0;
else reg_7c584cdd_u0<=reg_0ea303a6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2fda3f5d_u0<=1'h0;
else reg_2fda3f5d_u0<=reg_5421084c_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_46180292_u0<=1'h0;
else reg_46180292_u0<=reg_7fea3339_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3e132299_u0<=1'h0;
else reg_3e132299_u0<=reg_3bdd9bc2_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6b869f0a_u0<=1'h0;
else reg_6b869f0a_u0<=reg_5091952b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4f7f23f2_u0<=1'h0;
else reg_4f7f23f2_u0<=reg_5dc60849_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_133b2fb4_u0<=1'h0;
else reg_133b2fb4_u0<=reg_72251f10_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_64362ca6_u0<=1'h0;
else reg_64362ca6_u0<=reg_07fe52f5_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4ecc7e59_u0<=1'h0;
else reg_4ecc7e59_u0<=reg_2db318e2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3f4f33d9_u0<=1'h0;
else reg_3f4f33d9_u0<=reg_4d587466_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7399b70f_u0<=1'h0;
else reg_7399b70f_u0<=reg_6b869f0a_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_09c14556_u0<=1'h0;
else reg_09c14556_u0<=reg_5e91ea5a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_46180292_result_delayed_u0<=1'h0;
else reg_46180292_result_delayed_u0<=reg_46180292_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4e37ba53_result_delayed_u0<=1'h0;
else reg_4e37ba53_result_delayed_u0<=reg_4e37ba53_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_46e39e7c_u0<=1'h0;
else reg_46e39e7c_u0<=reg_40f72c06_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5aa3a23c_u0<=1'h0;
else reg_5aa3a23c_u0<=reg_4f7f23f2_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6a5362cc_u0<=1'h0;
else reg_6a5362cc_u0<=reg_2177b168_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6bfdef5c_u0<=1'h0;
else reg_6bfdef5c_u0<=reg_459701b4_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4f435be2_u0<=1'h0;
else reg_4f435be2_u0<=reg_12415e78_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_686a8c2c_result_delayed_u0<=1'h0;
else reg_686a8c2c_result_delayed_u0<=reg_686a8c2c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7136b992_u0<=1'h0;
else reg_7136b992_u0<=reg_05509604_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_30e39c45_u0<=1'h0;
else reg_30e39c45_u0<=reg_1d5b7d72_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2e5316fb_u0<=1'h0;
else reg_2e5316fb_u0<=reg_02899a41_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7f08dfa4_u0<=1'h0;
else reg_7f08dfa4_u0<=reg_56c7f61c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0bddd372_u0<=1'h0;
else reg_0bddd372_u0<=reg_5feeefb2_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_35cd15db_result_delayed_u0<=1'h0;
else reg_35cd15db_result_delayed_u0<=reg_35cd15db_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_39cf897d_u0<=1'h0;
else reg_39cf897d_u0<=reg_53cd0b25_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_42ddc26b_u0<=1'h0;
else reg_42ddc26b_u0<=reg_5c28119c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2cf5744d_u0<=1'h0;
else reg_2cf5744d_u0<=reg_39cf897d_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_03c03f7a_u0<=1'h0;
else reg_03c03f7a_u0<=reg_295e5824_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1941b9ff_u0<=1'h0;
else reg_1941b9ff_u0<=reg_658e74db_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3ddee161_u0<=1'h0;
else reg_3ddee161_u0<=reg_0a125ef3_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_215ed100_result_delayed_u0<=1'h0;
else reg_215ed100_result_delayed_u0<=reg_215ed100_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3ddee161_result_delayed_u0<=1'h0;
else reg_3ddee161_result_delayed_u0<=reg_3ddee161_u0;
end
assign or_u793_u0=and_delayed_u174|reg_09485a92_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_357fadb7_u0<=1'h0;
else reg_357fadb7_u0<=reg_6d8ffc20_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_02899a41_u0<=1'h0;
else reg_02899a41_u0<=reg_1b3d5a52_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2cf5703d_u0<=1'h0;
else reg_2cf5703d_u0<=reg_1941b9ff_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5e91ea5a_u0<=1'h0;
else reg_5e91ea5a_u0<=reg_6fa4028c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_133b2fb4_result_delayed_u0<=1'h0;
else reg_133b2fb4_result_delayed_u0<=reg_133b2fb4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3582bd53_u0<=1'h0;
else reg_3582bd53_u0<=reg_575abe47_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_33c9371a_u0<=1'h0;
else reg_33c9371a_u0<=reg_0bddd372_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7fea3339_u0<=1'h0;
else reg_7fea3339_u0<=reg_47f45fc0_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_328a525c_u0<=1'h0;
else reg_328a525c_u0<=reg_58641d44_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_38c2bc14_u0<=1'h0;
else reg_38c2bc14_u0<=reg_4d591d1c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0a55fe82_u0<=1'h0;
else reg_0a55fe82_u0<=reg_710aad0d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_357fadb7_result_delayed_u0<=1'h0;
else reg_357fadb7_result_delayed_u0<=reg_357fadb7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_50915049_u0<=1'h0;
else reg_50915049_u0<=reg_7ab59fff_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_742b90f1_u0<=1'h0;
else reg_742b90f1_u0<=reg_01f5f8bd_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_56c7f61c_u0<=1'h0;
else reg_56c7f61c_u0<=reg_2abca780_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_377e6fa5_u0<=1'h0;
else reg_377e6fa5_u0<=reg_7c7f2949_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_50915049_result_delayed_u0<=1'h0;
else reg_50915049_result_delayed_u0<=reg_50915049_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2cf5703d_result_delayed_u0<=1'h0;
else reg_2cf5703d_result_delayed_u0<=reg_2cf5703d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_42f8ea27_u0<=1'h0;
else reg_42f8ea27_u0<=reg_13f4d67d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7fea3339_result_delayed_u0<=1'h0;
else reg_7fea3339_result_delayed_u0<=reg_7fea3339_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0a125ef3_u0<=1'h0;
else reg_0a125ef3_u0<=reg_2a4e2976_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3ddee161_result_delayed_result_delayed_u0<=1'h0;
else reg_3ddee161_result_delayed_result_delayed_u0<=reg_3ddee161_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4f70c32f_result_delayed_u0<=1'h0;
else reg_4f70c32f_result_delayed_u0<=reg_4f70c32f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_67074bef_u0<=1'h0;
else reg_67074bef_u0<=reg_2e5316fb_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_53cd0b25_u0<=1'h0;
else reg_53cd0b25_u0<=reg_790c1f8e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4ecc7e59_result_delayed_u0<=1'h0;
else reg_4ecc7e59_result_delayed_u0<=reg_4ecc7e59_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_50915049_result_delayed_result_delayed_u0<=1'h0;
else reg_50915049_result_delayed_result_delayed_u0<=reg_50915049_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_47f45fc0_result_delayed_u0<=1'h0;
else reg_47f45fc0_result_delayed_u0<=reg_47f45fc0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_40f72c06_u0<=1'h0;
else reg_40f72c06_u0<=reg_0963c64e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7bbff74c_u0<=1'h0;
else reg_7bbff74c_u0<=reg_72076745_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3dda652e_u0<=1'h0;
else reg_3dda652e_u0<=reg_7d04d098_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3fc46730_u0<=1'h0;
else reg_3fc46730_u0<=reg_12fa7fcd_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7f74a383_u0<=1'h0;
else reg_7f74a383_u0<=reg_5b704959_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_42ddc26b_result_delayed_u0<=1'h0;
else reg_42ddc26b_result_delayed_u0<=reg_42ddc26b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4f6a4392_u0<=1'h0;
else reg_4f6a4392_u0<=reg_4b8c12d0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_331527ef_u0<=1'h0;
else reg_331527ef_u0<=reg_328a525c_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1e29aad3_u0<=1'h0;
else reg_1e29aad3_u0<=reg_3893a2cc_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3fd1972f_u0<=1'h0;
else reg_3fd1972f_u0<=reg_33d17fbe_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0ea303a6_u0<=1'h0;
else reg_0ea303a6_u0<=reg_382559bf_result_delayed_u0;
end
assign and_u2687_u0=and_u2682_u0&and_u2689_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4cade9aa_u0<=1'h0;
else reg_4cade9aa_u0<=reg_2defdc44_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6052ed5a_u0<=1'h0;
else reg_6052ed5a_u0<=reg_2892d198_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5421084c_result_delayed_u0<=1'h0;
else reg_5421084c_result_delayed_u0<=reg_5421084c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_20d8e0b0_result_delayed_u0<=1'h0;
else reg_20d8e0b0_result_delayed_u0<=reg_20d8e0b0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2892d198_u0<=1'h0;
else reg_2892d198_u0<=reg_7c584cdd_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_23e976e3_u0<=1'h0;
else reg_23e976e3_u0<=reg_6a5362cc_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_07fe52f5_u0<=1'h0;
else reg_07fe52f5_u0<=reg_377e6fa5_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7f74a383_result_delayed_u0<=1'h0;
else reg_7f74a383_result_delayed_u0<=reg_7f74a383_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_03bbbeb5_u0<=1'h0;
else reg_03bbbeb5_u0<=reg_41e078cd_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00a555b0_u0<=1'h0;
else reg_00a555b0_u0<=reg_3e2b8c33_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_16d553cc_u0<=1'h0;
else reg_16d553cc_u0<=reg_6ee35aab_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_45a48cbd_u0<=1'h0;
else reg_45a48cbd_u0<=reg_42ddc26b_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2cf5744d_result_delayed_u0<=1'h0;
else reg_2cf5744d_result_delayed_u0<=reg_2cf5744d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_459701b4_result_delayed_u0<=1'h0;
else reg_459701b4_result_delayed_u0<=reg_459701b4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3fd572c8_u0<=1'h0;
else reg_3fd572c8_u0<=reg_2cc01ca0_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_575abe47_u0<=1'h0;
else reg_575abe47_u0<=reg_74ed74eb_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_353a7c24_u0<=1'h0;
else reg_353a7c24_u0<=reg_3e561e48_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_58641d44_u0<=1'h0;
else reg_58641d44_u0<=reg_7ac1bb42_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6a5362cc_result_delayed_u0<=1'h0;
else reg_6a5362cc_result_delayed_u0<=reg_6a5362cc_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_25d144f5_u0<=1'h0;
else reg_25d144f5_u0<=reg_353a7c24_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6cdb19fe_u0<=1'h0;
else reg_6cdb19fe_u0<=reg_4497f4d9_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6fa4028c_u0<=1'h0;
else reg_6fa4028c_u0<=reg_6ca72548_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_41e078cd_u0<=1'h0;
else reg_41e078cd_u0<=reg_345a7803_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1fd68ee4_u0<=1'h0;
else reg_1fd68ee4_u0<=reg_133b2fb4_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7e0acb38_u0<=1'h0;
else reg_7e0acb38_u0<=reg_2cf5744d_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_72251f10_u0<=1'h0;
else reg_72251f10_u0<=reg_735e96ed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2cf5703d_result_delayed_result_delayed_u0<=1'h0;
else reg_2cf5703d_result_delayed_result_delayed_u0<=reg_2cf5703d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7c7f2949_u0<=1'h0;
else reg_7c7f2949_u0<=reg_0054d249_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2cc3d1f5_u0<=1'h0;
else reg_2cc3d1f5_u0<=reg_250a9f11_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_12fa7fcd_u0<=1'h0;
else reg_12fa7fcd_u0<=reg_571dd692_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2177b168_result_delayed_u0<=1'h0;
else reg_2177b168_result_delayed_u0<=reg_2177b168_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2abca780_u0<=1'h0;
else reg_2abca780_u0<=reg_4e9416d8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_71dddce1_u0<=1'h0;
else reg_71dddce1_u0<=reg_1d65b7da_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4d587466_u0<=1'h0;
else reg_4d587466_u0<=reg_0a55fe82_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_72076745_u0<=1'h0;
else reg_72076745_u0<=reg_607d9479_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6ff6deb2_u0<=1'h0;
else reg_6ff6deb2_u0<=reg_5fbaaa33_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3d9590d0_u0<=1'h0;
else reg_3d9590d0_u0<=reg_55043b64_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01f5f8bd_u0<=1'h0;
else reg_01f5f8bd_u0<=reg_62f7e6e1_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1a8e23c7_u0<=1'h0;
else reg_1a8e23c7_u0<=reg_0e5cbc7b_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7ab59fff_u0<=1'h0;
else reg_7ab59fff_u0<=reg_1d95898b_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4e37ba53_result_delayed_result_delayed_u0<=1'h0;
else reg_4e37ba53_result_delayed_result_delayed_u0<=reg_4e37ba53_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7bbff74c_result_delayed_u0<=1'h0;
else reg_7bbff74c_result_delayed_u0<=reg_7bbff74c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_77c337a8_result_delayed_u0<=1'h0;
else reg_77c337a8_result_delayed_u0<=reg_77c337a8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2892d198_result_delayed_u0<=1'h0;
else reg_2892d198_result_delayed_u0<=reg_2892d198_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6b869f0a_result_delayed_u0<=1'h0;
else reg_6b869f0a_result_delayed_u0<=reg_6b869f0a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2db318e2_u0<=1'h0;
else reg_2db318e2_u0<=reg_01347069_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_57c45696_u0<=1'h0;
else reg_57c45696_u0<=reg_2e407063_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_658e74db_u0<=1'h0;
else reg_658e74db_u0<=reg_38c2bc14_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_38c2bc14_result_delayed_u0<=1'h0;
else reg_38c2bc14_result_delayed_u0<=reg_38c2bc14_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4b8c12d0_u0<=1'h0;
else reg_4b8c12d0_u0<=reg_2e8ff2a2_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01347069_u0<=1'h0;
else reg_01347069_u0<=reg_63f53a08_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4e37ba53_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_4e37ba53_result_delayed_result_delayed_result_delayed_u0<=reg_4e37ba53_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_328a525c_result_delayed_u0<=1'h0;
else reg_328a525c_result_delayed_u0<=reg_328a525c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2cc3d1f5_result_delayed_u0<=1'h0;
else reg_2cc3d1f5_result_delayed_u0<=reg_2cc3d1f5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1c090d6c_u0<=1'h0;
else reg_1c090d6c_u0<=reg_46e39e7c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_33c9371a_result_delayed_u0<=1'h0;
else reg_33c9371a_result_delayed_u0<=reg_33c9371a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3851f050_result_delayed_u0<=1'h0;
else reg_3851f050_result_delayed_u0<=reg_3851f050_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2e8ff2a2_result_delayed_u0<=1'h0;
else reg_2e8ff2a2_result_delayed_u0<=reg_2e8ff2a2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0414817f_u0<=1'h0;
else reg_0414817f_u0<=reg_6bf27e46_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_185bb135_u0<=1'h0;
else reg_185bb135_u0<=reg_4e6c385a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1b3d5a52_u0<=1'h0;
else reg_1b3d5a52_u0<=reg_3e132299_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2c350944_u0<=1'h0;
else reg_2c350944_u0<=reg_7f74a383_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2af4ab86_u0<=1'h0;
else reg_2af4ab86_u0<=reg_53b43e36_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3113d461_u0<=1'h0;
else reg_3113d461_u0<=reg_77c337a8_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_295e5824_u0<=1'h0;
else reg_295e5824_u0<=reg_6cdb19fe_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_46180292_result_delayed_result_delayed_u0<=1'h0;
else reg_46180292_result_delayed_result_delayed_u0<=reg_46180292_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_38ae08a8_result_delayed_result_delayed_u0<=1'h0;
else reg_38ae08a8_result_delayed_result_delayed_u0<=reg_38ae08a8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5e62c71d_u0<=1'h0;
else reg_5e62c71d_u0<=reg_27aff15e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_44757003_result_delayed_u0<=1'h0;
else reg_44757003_result_delayed_u0<=reg_44757003_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7136b992_result_delayed_u0<=1'h0;
else reg_7136b992_result_delayed_u0<=reg_7136b992_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_53b43e36_u0<=1'h0;
else reg_53b43e36_u0<=reg_357fadb7_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_377e6fa5_result_delayed_u0<=1'h0;
else reg_377e6fa5_result_delayed_u0<=reg_377e6fa5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7ac1bb42_u0<=1'h0;
else reg_7ac1bb42_u0<=reg_6c3dc470_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7fd56e50_u0<=1'h0;
else reg_7fd56e50_u0<=reg_0b46a87d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_119a281f_u0<=1'h0;
else reg_119a281f_u0<=reg_2fda3f5d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_119a281f_result_delayed_u0<=1'h0;
else reg_119a281f_result_delayed_u0<=reg_119a281f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_030ef688_u0<=1'h0;
else reg_030ef688_u0<=reg_15ccc01d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_42ddc26b_result_delayed_result_delayed_u0<=1'h0;
else reg_42ddc26b_result_delayed_result_delayed_u0<=reg_42ddc26b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_13f4d67d_u0<=1'h0;
else reg_13f4d67d_u0<=reg_65138d26_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5fbaaa33_u0<=1'h0;
else reg_5fbaaa33_u0<=reg_398565f1_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_032d42a6_u0<=1'h0;
else reg_032d42a6_u0<=reg_4ba6c3eb_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5dc60849_u0<=1'h0;
else reg_5dc60849_u0<=reg_03bbbeb5_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_571dd692_u0<=1'h0;
else reg_571dd692_u0<=reg_1df705ad_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4ba6c3eb_result_delayed_u0<=1'h0;
else reg_4ba6c3eb_result_delayed_u0<=reg_4ba6c3eb_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_382559bf_u0<=1'h0;
else reg_382559bf_u0<=reg_072c9294_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_19da6841_u0<=1'h0;
else reg_19da6841_u0<=reg_5d8a9f60_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7d04d098_u0<=1'h0;
else reg_7d04d098_u0<=reg_2b8f21ae_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6ee35aab_result_delayed_u0<=1'h0;
else reg_6ee35aab_result_delayed_u0<=reg_6ee35aab_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7d04d098_result_delayed_u0<=1'h0;
else reg_7d04d098_result_delayed_u0<=reg_7d04d098_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0ef27753_u0<=1'h0;
else reg_0ef27753_u0<=reg_38ae08a8_result_delayed_result_delayed_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6ff6deb2_result_delayed_u0<=1'h0;
else reg_6ff6deb2_result_delayed_u0<=reg_6ff6deb2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1d5b7d72_result_delayed_u0<=1'h0;
else reg_1d5b7d72_result_delayed_u0<=reg_1d5b7d72_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2defdc44_u0<=1'h0;
else reg_2defdc44_u0<=reg_4a16e8d3_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5bba6fd9_result_delayed_u0<=1'h0;
else reg_5bba6fd9_result_delayed_u0<=reg_5bba6fd9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01f5f8bd_result_delayed_u0<=1'h0;
else reg_01f5f8bd_result_delayed_u0<=reg_01f5f8bd_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6d8ffc20_u0<=1'h0;
else reg_6d8ffc20_u0<=reg_11bf5a5d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6cdb19fe_result_delayed_u0<=1'h0;
else reg_6cdb19fe_result_delayed_u0<=reg_6cdb19fe_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7f74a383_result_delayed_result_delayed_u0<=1'h0;
else reg_7f74a383_result_delayed_result_delayed_u0<=reg_7f74a383_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_735e96ed_u0<=1'h0;
else reg_735e96ed_u0<=reg_44757003_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6bf27e46_u0<=1'h0;
else reg_6bf27e46_u0<=reg_5aa3a23c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5c28119c_u0<=1'h0;
else reg_5c28119c_u0<=reg_3dda652e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_07aa93c1_result_delayed_u0<=1'h0;
else reg_07aa93c1_result_delayed_u0<=reg_07aa93c1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_072c9294_u0<=1'h0;
else reg_072c9294_u0<=reg_3fd1972f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5091952b_u0<=1'h0;
else reg_5091952b_u0<=reg_2be729d4_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7ce31523_u0<=1'h0;
else reg_7ce31523_u0<=reg_2d137930_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_25d144f5_result_delayed_u0<=1'h0;
else reg_25d144f5_result_delayed_u0<=reg_25d144f5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_12415e78_result_delayed_u0<=1'h0;
else reg_12415e78_result_delayed_u0<=reg_12415e78_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_35cd15db_result_delayed_result_delayed_u0<=1'h0;
else reg_35cd15db_result_delayed_result_delayed_u0<=reg_35cd15db_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_40f72c06_result_delayed_u0<=1'h0;
else reg_40f72c06_result_delayed_u0<=reg_40f72c06_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3e561e48_result_delayed_u0<=1'h0;
else reg_3e561e48_result_delayed_u0<=reg_3e561e48_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_57c45696_result_delayed_u0<=1'h0;
else reg_57c45696_result_delayed_u0<=reg_57c45696_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6a6f9fa5_u0<=1'h0;
else reg_6a6f9fa5_u0<=reg_33c9371a_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7c87d14d_u0<=1'h0;
else reg_7c87d14d_u0<=reg_7399b70f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0ef27753_result_delayed_u0<=1'h0;
else reg_0ef27753_result_delayed_u0<=reg_0ef27753_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00a555b0_result_delayed_u0<=1'h0;
else reg_00a555b0_result_delayed_u0<=reg_00a555b0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1941b9ff_result_delayed_u0<=1'h0;
else reg_1941b9ff_result_delayed_u0<=reg_1941b9ff_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_28b4d165_u0<=1'h0;
else reg_28b4d165_u0<=reg_3fd572c8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_15ccc01d_u0<=1'h0;
else reg_15ccc01d_u0<=reg_023bffd6_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2cc3d1f5_result_delayed_result_delayed_u0<=1'h0;
else reg_2cc3d1f5_result_delayed_result_delayed_u0<=reg_2cc3d1f5_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_09c14556_result_delayed_u0<=1'h0;
else reg_09c14556_result_delayed_u0<=reg_09c14556_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_32854b5c_u0<=1'h0;
else reg_32854b5c_u0<=reg_2a22ac7d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6134ccef_u0<=1'h0;
else reg_6134ccef_u0<=reg_79022b5e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7572dd7f_result_delayed_u0<=1'h0;
else reg_7572dd7f_result_delayed_u0<=reg_7572dd7f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_30e39c45_result_delayed_u0<=1'h0;
else reg_30e39c45_result_delayed_u0<=reg_30e39c45_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6ed66f32_u0<=1'h0;
else reg_6ed66f32_u0<=reg_4cf0ecf8_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_78342dd1_u0<=1'h0;
else reg_78342dd1_u0<=reg_20d8e0b0_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0f9d1678_u0<=1'h0;
else reg_0f9d1678_u0<=reg_3851f050_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0414817f_result_delayed_u0<=1'h0;
else reg_0414817f_result_delayed_u0<=reg_0414817f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4f852262_u0<=1'h0;
else reg_4f852262_u0<=reg_0f9d1678_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_023bffd6_u0<=1'h0;
else reg_023bffd6_u0<=reg_7572dd7f_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_596f7c82_u0<=1'h0;
else reg_596f7c82_u0<=reg_1f57f175_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6ca72548_u0<=1'h0;
else reg_6ca72548_u0<=reg_4cade9aa_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1fd68ee4_result_delayed_u0<=1'h0;
else reg_1fd68ee4_result_delayed_u0<=reg_1fd68ee4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_07fe52f5_result_delayed_u0<=1'h0;
else reg_07fe52f5_result_delayed_u0<=reg_07fe52f5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_16d553cc_result_delayed_u0<=1'h0;
else reg_16d553cc_result_delayed_u0<=reg_16d553cc_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1b102eec_u0<=1'h0;
else reg_1b102eec_u0<=reg_71dddce1_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_63f53a08_u0<=1'h0;
else reg_63f53a08_u0<=reg_35cd15db_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_38ae08a8_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_38ae08a8_result_delayed_result_delayed_result_delayed_u0<=reg_38ae08a8_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4cade9aa_result_delayed_u0<=1'h0;
else reg_4cade9aa_result_delayed_u0<=reg_4cade9aa_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_795d0757_u0<=1'h0;
else reg_795d0757_u0<=reg_6134ccef_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_44757003_result_delayed_result_delayed_u0<=1'h0;
else reg_44757003_result_delayed_result_delayed_u0<=reg_44757003_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_751aa708_u0<=1'h0;
else reg_751aa708_u0<=reg_3113d461_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1479ea6c_u0<=1'h0;
else reg_1479ea6c_u0<=reg_45a48cbd_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_33c9371a_result_delayed_result_delayed_u0<=1'h0;
else reg_33c9371a_result_delayed_result_delayed_u0<=reg_33c9371a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3e2b8c33_u0<=1'h0;
else reg_3e2b8c33_u0<=reg_7bbff74c_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2af4ab86_result_delayed_u0<=1'h0;
else reg_2af4ab86_result_delayed_u0<=reg_2af4ab86_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1941b9ff_result_delayed_result_delayed_u0<=1'h0;
else reg_1941b9ff_result_delayed_result_delayed_u0<=reg_1941b9ff_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_250a9f11_u0<=1'h0;
else reg_250a9f11_u0<=reg_4ecc7e59_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7b11510d_u0<=1'h0;
else reg_7b11510d_u0<=reg_686a8c2c_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4497f4d9_result_delayed_u0<=1'h0;
else reg_4497f4d9_result_delayed_u0<=reg_4497f4d9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_39cf897d_result_delayed_u0<=1'h0;
else reg_39cf897d_result_delayed_u0<=reg_39cf897d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0054d249_u0<=1'h0;
else reg_0054d249_u0<=reg_6aa4982f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_74ed74eb_result_delayed_u0<=1'h0;
else reg_74ed74eb_result_delayed_u0<=reg_74ed74eb_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2b8f21ae_u0<=1'h0;
else reg_2b8f21ae_u0<=reg_2c350944_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1f57f175_u0<=1'h0;
else reg_1f57f175_u0<=reg_43fabda0_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_28b4d165_result_delayed_u0<=1'h0;
else reg_28b4d165_result_delayed_u0<=reg_28b4d165_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2e407063_u0<=1'h0;
else reg_2e407063_u0<=reg_6761984a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0e5cbc7b_u0<=1'h0;
else reg_0e5cbc7b_u0<=reg_3fc46730_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5b704959_u0<=1'h0;
else reg_5b704959_u0<=reg_7ce31523_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4f7f23f2_result_delayed_u0<=1'h0;
else reg_4f7f23f2_result_delayed_u0<=reg_4f7f23f2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6ed66f32_result_delayed_u0<=1'h0;
else reg_6ed66f32_result_delayed_u0<=reg_6ed66f32_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_357fadb7_result_delayed_result_delayed_u0<=1'h0;
else reg_357fadb7_result_delayed_result_delayed_u0<=reg_357fadb7_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_03bbbeb5_result_delayed_u0<=1'h0;
else reg_03bbbeb5_result_delayed_u0<=reg_03bbbeb5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2be729d4_u0<=1'h0;
else reg_2be729d4_u0<=reg_14905eff_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_63f53a08_result_delayed_u0<=1'h0;
else reg_63f53a08_result_delayed_u0<=reg_63f53a08_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4e6c385a_u0<=1'h0;
else reg_4e6c385a_u0<=reg_23e976e3_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0bddd372_result_delayed_u0<=1'h0;
else reg_0bddd372_result_delayed_u0<=reg_0bddd372_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2cf5744d_result_delayed_result_delayed_u0<=1'h0;
else reg_2cf5744d_result_delayed_result_delayed_u0<=reg_2cf5744d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0576bf35_u0<=1'h0;
else reg_0576bf35_u0<=reg_3cf3ff64_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_33d17fbe_result_delayed_u0<=1'h0;
else reg_33d17fbe_result_delayed_u0<=reg_33d17fbe_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_14095c65_result_delayed_u0<=1'h0;
else reg_14095c65_result_delayed_u0<=reg_14095c65_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_46e39e7c_result_delayed_u0<=1'h0;
else reg_46e39e7c_result_delayed_u0<=reg_46e39e7c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2cc01ca0_result_delayed_u0<=1'h0;
else reg_2cc01ca0_result_delayed_u0<=reg_2cc01ca0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7ac1bb42_result_delayed_u0<=1'h0;
else reg_7ac1bb42_result_delayed_u0<=reg_7ac1bb42_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4d587466_result_delayed_u0<=1'h0;
else reg_4d587466_result_delayed_u0<=reg_4d587466_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_45a48cbd_result_delayed_u0<=1'h0;
else reg_45a48cbd_result_delayed_u0<=reg_45a48cbd_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2cfcc2a4_u0<=1'h0;
else reg_2cfcc2a4_u0<=reg_7fd56e50_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_43fabda0_u0<=1'h0;
else reg_43fabda0_u0<=reg_1a8e23c7_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_79022b5e_u0<=1'h0;
else reg_79022b5e_u0<=reg_738977bb_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3fc46730_result_delayed_u0<=1'h0;
else reg_3fc46730_result_delayed_u0<=reg_3fc46730_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_35cd15db_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_35cd15db_result_delayed_result_delayed_result_delayed_u0<=reg_35cd15db_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2a22ac7d_u0<=1'h0;
else reg_2a22ac7d_u0<=reg_119a281f_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3893a2cc_u0<=1'h0;
else reg_3893a2cc_u0<=reg_2bfc93f9_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_55043b64_u0<=1'h0;
else reg_55043b64_u0<=reg_30e39c45_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6134ccef_result_delayed_u0<=1'h0;
else reg_6134ccef_result_delayed_u0<=reg_6134ccef_u0;
end
assign and_u2688_u0=and_u2683_u0&and_u2689_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_58980aff_u0<=1'h0;
else reg_58980aff_u0<=reg_4f70c32f_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3156ef3e_u0<=1'h0;
else reg_3156ef3e_u0<=reg_25d144f5_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5feeefb2_result_delayed_u0<=1'h0;
else reg_5feeefb2_result_delayed_u0<=reg_5feeefb2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_14905eff_u0<=1'h0;
else reg_14905eff_u0<=reg_0b346188_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_03bbbeb5_result_delayed_result_delayed_u0<=1'h0;
else reg_03bbbeb5_result_delayed_result_delayed_u0<=reg_03bbbeb5_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_07fe52f5_result_delayed_result_delayed_u0<=1'h0;
else reg_07fe52f5_result_delayed_result_delayed_u0<=reg_07fe52f5_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0576bf35_result_delayed_u0<=1'h0;
else reg_0576bf35_result_delayed_u0<=reg_0576bf35_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_30e39c45_result_delayed_result_delayed_u0<=1'h0;
else reg_30e39c45_result_delayed_result_delayed_u0<=reg_30e39c45_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3843f63d_u0<=1'h0;
else reg_3843f63d_u0<=reg_032d42a6_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01f5f8bd_result_delayed_result_delayed_u0<=1'h0;
else reg_01f5f8bd_result_delayed_result_delayed_u0<=reg_01f5f8bd_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2be729d4_result_delayed_u0<=1'h0;
else reg_2be729d4_result_delayed_u0<=reg_2be729d4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_79022b5e_result_delayed_u0<=1'h0;
else reg_79022b5e_result_delayed_u0<=reg_79022b5e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_23e976e3_result_delayed_u0<=1'h0;
else reg_23e976e3_result_delayed_u0<=reg_23e976e3_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_790c1f8e_u0<=1'h0;
else reg_790c1f8e_u0<=reg_751aa708_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_47f45fc0_result_delayed_result_delayed_u0<=1'h0;
else reg_47f45fc0_result_delayed_result_delayed_u0<=reg_47f45fc0_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_217203f5_u0<=1'h0;
else reg_217203f5_u0<=reg_67074bef_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6aa4982f_u0<=1'h0;
else reg_6aa4982f_u0<=reg_3843f63d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_16d553cc_result_delayed_result_delayed_u0<=1'h0;
else reg_16d553cc_result_delayed_result_delayed_u0<=reg_16d553cc_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_795d0757_result_delayed_u0<=1'h0;
else reg_795d0757_result_delayed_u0<=reg_795d0757_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2cf5744d_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_2cf5744d_result_delayed_result_delayed_result_delayed_u0<=reg_2cf5744d_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4f70c32f_result_delayed_result_delayed_u0<=1'h0;
else reg_4f70c32f_result_delayed_result_delayed_u0<=reg_4f70c32f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2e5316fb_result_delayed_u0<=1'h0;
else reg_2e5316fb_result_delayed_u0<=reg_2e5316fb_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_04fc925c_u0<=1'h0;
else reg_04fc925c_u0<=reg_795d0757_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_62f7e6e1_result_delayed_u0<=1'h0;
else reg_62f7e6e1_result_delayed_u0<=reg_62f7e6e1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_710aad0d_result_delayed_u0<=1'h0;
else reg_710aad0d_result_delayed_u0<=reg_710aad0d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_32854b5c_result_delayed_u0<=1'h0;
else reg_32854b5c_result_delayed_u0<=reg_32854b5c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1d95898b_result_delayed_u0<=1'h0;
else reg_1d95898b_result_delayed_u0<=reg_1d95898b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_25d144f5_result_delayed_result_delayed_u0<=1'h0;
else reg_25d144f5_result_delayed_result_delayed_u0<=reg_25d144f5_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_686a8c2c_result_delayed_result_delayed_u0<=1'h0;
else reg_686a8c2c_result_delayed_result_delayed_u0<=reg_686a8c2c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_058dcb20_u0<=1'h0;
else reg_058dcb20_u0<=reg_46180292_result_delayed_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5bba6fd9_result_delayed_result_delayed_u0<=1'h0;
else reg_5bba6fd9_result_delayed_result_delayed_u0<=reg_5bba6fd9_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_43fabda0_result_delayed_u0<=1'h0;
else reg_43fabda0_result_delayed_u0<=reg_43fabda0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4f70c32f_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_4f70c32f_result_delayed_result_delayed_result_delayed_u0<=reg_4f70c32f_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5574bbc5_u0<=1'h0;
else reg_5574bbc5_u0<=reg_75d7ab69_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_607d9479_result_delayed_u0<=1'h0;
else reg_607d9479_result_delayed_u0<=reg_607d9479_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3fd1972f_result_delayed_u0<=1'h0;
else reg_3fd1972f_result_delayed_u0<=reg_3fd1972f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_38ae08a8_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_38ae08a8_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_38ae08a8_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6c3dc470_result_delayed_u0<=1'h0;
else reg_6c3dc470_result_delayed_u0<=reg_6c3dc470_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0b346188_u0<=1'h0;
else reg_0b346188_u0<=reg_1b102eec_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_38ae08a8_result_delayed_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_38ae08a8_result_delayed_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_38ae08a8_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7572dd7f_result_delayed_result_delayed_u0<=1'h0;
else reg_7572dd7f_result_delayed_result_delayed_u0<=reg_7572dd7f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_75d7ab69_u0<=1'h0;
else reg_75d7ab69_u0<=reg_1eed982d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1d65b7da_u0<=1'h0;
else reg_1d65b7da_u0<=reg_2cbb2cce_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1eed982d_u0<=1'h0;
else reg_1eed982d_u0<=reg_185bb135_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1479ea6c_result_delayed_u0<=1'h0;
else reg_1479ea6c_result_delayed_u0<=reg_1479ea6c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_42f8ea27_result_delayed_u0<=1'h0;
else reg_42f8ea27_result_delayed_u0<=reg_42f8ea27_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4a16e8d3_u0<=1'h0;
else reg_4a16e8d3_u0<=reg_7b11510d_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2cf5744d_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_2cf5744d_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_2cf5744d_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2be729d4_result_delayed_result_delayed_u0<=1'h0;
else reg_2be729d4_result_delayed_result_delayed_u0<=reg_2be729d4_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3893a2cc_result_delayed_u0<=1'h0;
else reg_3893a2cc_result_delayed_u0<=reg_3893a2cc_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5aa3a23c_result_delayed_u0<=1'h0;
else reg_5aa3a23c_result_delayed_u0<=reg_5aa3a23c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_051b0973_result_delayed_u0<=1'h0;
else reg_051b0973_result_delayed_u0<=reg_051b0973_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_331527ef_result_delayed_u0<=1'h0;
else reg_331527ef_result_delayed_u0<=reg_331527ef_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01347069_result_delayed_u0<=1'h0;
else reg_01347069_result_delayed_u0<=reg_01347069_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3fd572c8_result_delayed_u0<=1'h0;
else reg_3fd572c8_result_delayed_u0<=reg_3fd572c8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_20d8e0b0_result_delayed_result_delayed_u0<=1'h0;
else reg_20d8e0b0_result_delayed_result_delayed_u0<=reg_20d8e0b0_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_12415e78_result_delayed_result_delayed_u0<=1'h0;
else reg_12415e78_result_delayed_result_delayed_u0<=reg_12415e78_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6d8ffc20_result_delayed_u0<=1'h0;
else reg_6d8ffc20_result_delayed_u0<=reg_6d8ffc20_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_738977bb_result_delayed_u0<=1'h0;
else reg_738977bb_result_delayed_u0<=reg_738977bb_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6ff6deb2_result_delayed_result_delayed_u0<=1'h0;
else reg_6ff6deb2_result_delayed_result_delayed_u0<=reg_6ff6deb2_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_658e74db_result_delayed_u0<=1'h0;
else reg_658e74db_result_delayed_u0<=reg_658e74db_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5d8a9f60_u0<=1'h0;
else reg_5d8a9f60_u0<=reg_331527ef_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_30e39c45_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_30e39c45_result_delayed_result_delayed_result_delayed_u0<=reg_30e39c45_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_023bffd6_result_delayed_u0<=1'h0;
else reg_023bffd6_result_delayed_u0<=reg_023bffd6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4e9416d8_result_delayed_u0<=1'h0;
else reg_4e9416d8_result_delayed_u0<=reg_4e9416d8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_27aff15e_u0<=1'h0;
else reg_27aff15e_u0<=reg_051b0973_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_331527ef_result_delayed_result_delayed_u0<=1'h0;
else reg_331527ef_result_delayed_result_delayed_u0<=reg_331527ef_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_30e39c45_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_30e39c45_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_30e39c45_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_353a7c24_result_delayed_u0<=1'h0;
else reg_353a7c24_result_delayed_u0<=reg_353a7c24_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5d8a9f60_result_delayed_u0<=1'h0;
else reg_5d8a9f60_result_delayed_u0<=reg_5d8a9f60_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2892d198_result_delayed_result_delayed_u0<=1'h0;
else reg_2892d198_result_delayed_result_delayed_u0<=reg_2892d198_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2cbb2cce_result_delayed_u0<=1'h0;
else reg_2cbb2cce_result_delayed_u0<=reg_2cbb2cce_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7136b992_result_delayed_result_delayed_u0<=1'h0;
else reg_7136b992_result_delayed_result_delayed_u0<=reg_7136b992_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_133b2fb4_result_delayed_result_delayed_u0<=1'h0;
else reg_133b2fb4_result_delayed_result_delayed_u0<=reg_133b2fb4_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0a55fe82_result_delayed_u0<=1'h0;
else reg_0a55fe82_result_delayed_u0<=reg_0a55fe82_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2892d198_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_2892d198_result_delayed_result_delayed_result_delayed_u0<=reg_2892d198_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7b11510d_result_delayed_u0<=1'h0;
else reg_7b11510d_result_delayed_u0<=reg_7b11510d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_795d0757_result_delayed_result_delayed_u0<=1'h0;
else reg_795d0757_result_delayed_result_delayed_u0<=reg_795d0757_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0e5cbc7b_result_delayed_u0<=1'h0;
else reg_0e5cbc7b_result_delayed_u0<=reg_0e5cbc7b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5421084c_result_delayed_result_delayed_u0<=1'h0;
else reg_5421084c_result_delayed_result_delayed_u0<=reg_5421084c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7c584cdd_result_delayed_u0<=1'h0;
else reg_7c584cdd_result_delayed_u0<=reg_7c584cdd_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_571dd692_result_delayed_u0<=1'h0;
else reg_571dd692_result_delayed_u0<=reg_571dd692_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_575abe47_result_delayed_u0<=1'h0;
else reg_575abe47_result_delayed_u0<=reg_575abe47_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_12fa7fcd_result_delayed_u0<=1'h0;
else reg_12fa7fcd_result_delayed_u0<=reg_12fa7fcd_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_331527ef_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_331527ef_result_delayed_result_delayed_result_delayed_u0<=reg_331527ef_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_38ae08a8_result_delayed_result_delayed_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_38ae08a8_result_delayed_result_delayed_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_38ae08a8_result_delayed_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_658e74db_result_delayed_result_delayed_u0<=1'h0;
else reg_658e74db_result_delayed_result_delayed_u0<=reg_658e74db_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6761984a_u0<=1'h0;
else reg_6761984a_u0<=reg_0ef27753_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0963c64e_u0<=1'h0;
else reg_0963c64e_u0<=reg_57c45696_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3f4f33d9_result_delayed_u0<=1'h0;
else reg_3f4f33d9_result_delayed_u0<=reg_3f4f33d9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_751aa708_result_delayed_u0<=1'h0;
else reg_751aa708_result_delayed_u0<=reg_751aa708_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4ecc7e59_result_delayed_result_delayed_u0<=1'h0;
else reg_4ecc7e59_result_delayed_result_delayed_u0<=reg_4ecc7e59_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2a4e2976_u0<=1'h0;
else reg_2a4e2976_u0<=reg_31f2b9fa_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0b46a87d_u0<=1'h0;
else reg_0b46a87d_u0<=reg_6ff6deb2_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1eed982d_result_delayed_u0<=1'h0;
else reg_1eed982d_result_delayed_u0<=reg_1eed982d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6ed66f32_result_delayed_result_delayed_u0<=1'h0;
else reg_6ed66f32_result_delayed_result_delayed_u0<=reg_6ed66f32_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3113d461_result_delayed_u0<=1'h0;
else reg_3113d461_result_delayed_u0<=reg_3113d461_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3851f050_result_delayed_result_delayed_u0<=1'h0;
else reg_3851f050_result_delayed_result_delayed_u0<=reg_3851f050_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_67074bef_result_delayed_u0<=1'h0;
else reg_67074bef_result_delayed_u0<=reg_67074bef_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5b704959_result_delayed_u0<=1'h0;
else reg_5b704959_result_delayed_u0<=reg_5b704959_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_05509604_u0<=1'h0;
else reg_05509604_u0<=reg_1479ea6c_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3582bd53_result_delayed_u0<=1'h0;
else reg_3582bd53_result_delayed_u0<=reg_3582bd53_u0;
end
assign or_u794_u0=and_u2687_u0|and_u2686_u0;
assign mux_u270=(and_u2687_u0)?1'h1:1'h0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_46180292_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_46180292_result_delayed_result_delayed_result_delayed_u0<=reg_46180292_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2e5316fb_result_delayed_result_delayed_u0<=1'h0;
else reg_2e5316fb_result_delayed_result_delayed_u0<=reg_2e5316fb_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_46180292_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_46180292_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_46180292_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1b102eec_result_delayed_u0<=1'h0;
else reg_1b102eec_result_delayed_u0<=reg_1b102eec_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_39cf897d_result_delayed_result_delayed_u0<=1'h0;
else reg_39cf897d_result_delayed_result_delayed_u0<=reg_39cf897d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_459701b4_result_delayed_result_delayed_u0<=1'h0;
else reg_459701b4_result_delayed_result_delayed_u0<=reg_459701b4_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6ff6deb2_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_6ff6deb2_result_delayed_result_delayed_result_delayed_u0<=reg_6ff6deb2_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7d04d098_result_delayed_result_delayed_u0<=1'h0;
else reg_7d04d098_result_delayed_result_delayed_u0<=reg_7d04d098_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_58980aff_result_delayed_u0<=1'h0;
else reg_58980aff_result_delayed_u0<=reg_58980aff_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7399b70f_result_delayed_u0<=1'h0;
else reg_7399b70f_result_delayed_u0<=reg_7399b70f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4ba6c3eb_result_delayed_result_delayed_u0<=1'h0;
else reg_4ba6c3eb_result_delayed_result_delayed_u0<=reg_4ba6c3eb_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3bdd9bc2_result_delayed_u0<=1'h0;
else reg_3bdd9bc2_result_delayed_u0<=reg_3bdd9bc2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2a4e2976_result_delayed_u0<=1'h0;
else reg_2a4e2976_result_delayed_u0<=reg_2a4e2976_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_382559bf_result_delayed_u0<=1'h0;
else reg_382559bf_result_delayed_u0<=reg_382559bf_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7fea3339_result_delayed_result_delayed_u0<=1'h0;
else reg_7fea3339_result_delayed_result_delayed_u0<=reg_7fea3339_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_32854b5c_result_delayed_result_delayed_u0<=1'h0;
else reg_32854b5c_result_delayed_result_delayed_u0<=reg_32854b5c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_75d7ab69_result_delayed_u0<=1'h0;
else reg_75d7ab69_result_delayed_u0<=reg_75d7ab69_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4497f4d9_result_delayed_result_delayed_u0<=1'h0;
else reg_4497f4d9_result_delayed_result_delayed_u0<=reg_4497f4d9_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4f435be2_result_delayed_u0<=1'h0;
else reg_4f435be2_result_delayed_u0<=reg_4f435be2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0f9d1678_result_delayed_u0<=1'h0;
else reg_0f9d1678_result_delayed_u0<=reg_0f9d1678_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7fd56e50_result_delayed_u0<=1'h0;
else reg_7fd56e50_result_delayed_u0<=reg_7fd56e50_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3e132299_result_delayed_u0<=1'h0;
else reg_3e132299_result_delayed_u0<=reg_3e132299_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2e5316fb_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_2e5316fb_result_delayed_result_delayed_result_delayed_u0<=reg_2e5316fb_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_098c01f7_result_delayed_u0<=1'h0;
else reg_098c01f7_result_delayed_u0<=reg_098c01f7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_032d42a6_result_delayed_u0<=1'h0;
else reg_032d42a6_result_delayed_u0<=reg_032d42a6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_65138d26_result_delayed_u0<=1'h0;
else reg_65138d26_result_delayed_u0<=reg_65138d26_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_57c45696_result_delayed_result_delayed_u0<=1'h0;
else reg_57c45696_result_delayed_result_delayed_u0<=reg_57c45696_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_742b90f1_result_delayed_u0<=1'h0;
else reg_742b90f1_result_delayed_u0<=reg_742b90f1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_78342dd1_result_delayed_u0<=1'h0;
else reg_78342dd1_result_delayed_u0<=reg_78342dd1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2bfc93f9_result_delayed_u0<=1'h0;
else reg_2bfc93f9_result_delayed_u0<=reg_2bfc93f9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6b869f0a_result_delayed_result_delayed_u0<=1'h0;
else reg_6b869f0a_result_delayed_result_delayed_u0<=reg_6b869f0a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0576bf35_result_delayed_result_delayed_u0<=1'h0;
else reg_0576bf35_result_delayed_result_delayed_u0<=reg_0576bf35_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0576bf35_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_0576bf35_result_delayed_result_delayed_result_delayed_u0<=reg_0576bf35_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7c7f2949_result_delayed_u0<=1'h0;
else reg_7c7f2949_result_delayed_u0<=reg_7c7f2949_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3cf3ff64_u0<=1'h0;
else reg_3cf3ff64_u0<=reg_07aa93c1_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_185bb135_result_delayed_u0<=1'h0;
else reg_185bb135_result_delayed_u0<=reg_185bb135_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7b11510d_result_delayed_result_delayed_u0<=1'h0;
else reg_7b11510d_result_delayed_result_delayed_u0<=reg_7b11510d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3bdd9bc2_result_delayed_result_delayed_u0<=1'h0;
else reg_3bdd9bc2_result_delayed_result_delayed_u0<=reg_3bdd9bc2_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1d65b7da_result_delayed_u0<=1'h0;
else reg_1d65b7da_result_delayed_u0<=reg_1d65b7da_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_398565f1_result_delayed_u0<=1'h0;
else reg_398565f1_result_delayed_u0<=reg_398565f1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6ca72548_result_delayed_u0<=1'h0;
else reg_6ca72548_result_delayed_u0<=reg_6ca72548_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_345a7803_result_delayed_u0<=1'h0;
else reg_345a7803_result_delayed_u0<=reg_345a7803_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5d8a9f60_result_delayed_result_delayed_u0<=1'h0;
else reg_5d8a9f60_result_delayed_result_delayed_u0<=reg_5d8a9f60_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_571dd692_result_delayed_result_delayed_u0<=1'h0;
else reg_571dd692_result_delayed_result_delayed_u0<=reg_571dd692_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_328a525c_result_delayed_result_delayed_u0<=1'h0;
else reg_328a525c_result_delayed_result_delayed_u0<=reg_328a525c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0a125ef3_result_delayed_u0<=1'h0;
else reg_0a125ef3_result_delayed_u0<=reg_0a125ef3_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3cf3ff64_result_delayed_u0<=1'h0;
else reg_3cf3ff64_result_delayed_u0<=reg_3cf3ff64_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4b4698ef_u0<=1'h0;
else reg_4b4698ef_u0<=reg_217203f5_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_07aa93c1_result_delayed_result_delayed_u0<=1'h0;
else reg_07aa93c1_result_delayed_result_delayed_u0<=reg_07aa93c1_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0e5cbc7b_result_delayed_result_delayed_u0<=1'h0;
else reg_0e5cbc7b_result_delayed_result_delayed_u0<=reg_0e5cbc7b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_14905eff_result_delayed_u0<=1'h0;
else reg_14905eff_result_delayed_u0<=reg_14905eff_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_051b0973_result_delayed_result_delayed_u0<=1'h0;
else reg_051b0973_result_delayed_result_delayed_u0<=reg_051b0973_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1df705ad_result_delayed_u0<=1'h0;
else reg_1df705ad_result_delayed_u0<=reg_1df705ad_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3dda652e_result_delayed_u0<=1'h0;
else reg_3dda652e_result_delayed_u0<=reg_3dda652e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2fda3f5d_result_delayed_u0<=1'h0;
else reg_2fda3f5d_result_delayed_u0<=reg_2fda3f5d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1479ea6c_result_delayed_result_delayed_u0<=1'h0;
else reg_1479ea6c_result_delayed_result_delayed_u0<=reg_1479ea6c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_217203f5_result_delayed_u0<=1'h0;
else reg_217203f5_result_delayed_u0<=reg_217203f5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1d95898b_result_delayed_result_delayed_u0<=1'h0;
else reg_1d95898b_result_delayed_result_delayed_u0<=reg_1d95898b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2a22ac7d_result_delayed_u0<=1'h0;
else reg_2a22ac7d_result_delayed_u0<=reg_2a22ac7d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2f3b2083_u0<=1'h0;
else reg_2f3b2083_u0<=reg_3582bd53_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_31f2b9fa_result_delayed_u0<=1'h0;
else reg_31f2b9fa_result_delayed_u0<=reg_31f2b9fa_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_119a281f_result_delayed_result_delayed_u0<=1'h0;
else reg_119a281f_result_delayed_result_delayed_u0<=reg_119a281f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_43fabda0_result_delayed_result_delayed_u0<=1'h0;
else reg_43fabda0_result_delayed_result_delayed_u0<=reg_43fabda0_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_31f2b9fa_result_delayed_result_delayed_u0<=1'h0;
else reg_31f2b9fa_result_delayed_result_delayed_u0<=reg_31f2b9fa_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_795d0757_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_795d0757_result_delayed_result_delayed_result_delayed_u0<=reg_795d0757_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6134ccef_result_delayed_result_delayed_u0<=1'h0;
else reg_6134ccef_result_delayed_result_delayed_u0<=reg_6134ccef_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_77c337a8_result_delayed_result_delayed_u0<=1'h0;
else reg_77c337a8_result_delayed_result_delayed_u0<=reg_77c337a8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_71dddce1_result_delayed_u0<=1'h0;
else reg_71dddce1_result_delayed_u0<=reg_71dddce1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2f3b2083_result_delayed_u0<=1'h0;
else reg_2f3b2083_result_delayed_u0<=reg_2f3b2083_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7ce31523_result_delayed_u0<=1'h0;
else reg_7ce31523_result_delayed_u0<=reg_7ce31523_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_459701b4_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_459701b4_result_delayed_result_delayed_result_delayed_u0<=reg_459701b4_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_09485a92_u0<=1'h0;
else reg_09485a92_u0<=reg_7c87d14d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3843f63d_result_delayed_u0<=1'h0;
else reg_3843f63d_result_delayed_u0<=reg_3843f63d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0ef27753_result_delayed_result_delayed_u0<=1'h0;
else reg_0ef27753_result_delayed_result_delayed_u0<=reg_0ef27753_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_23c003c5_result_delayed_u0<=1'h0;
else reg_23c003c5_result_delayed_u0<=reg_23c003c5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4f70c32f_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_4f70c32f_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_4f70c32f_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2cc01ca0_result_delayed_result_delayed_u0<=1'h0;
else reg_2cc01ca0_result_delayed_result_delayed_u0<=reg_2cc01ca0_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3582bd53_result_delayed_result_delayed_u0<=1'h0;
else reg_3582bd53_result_delayed_result_delayed_u0<=reg_3582bd53_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1a8e23c7_result_delayed_u0<=1'h0;
else reg_1a8e23c7_result_delayed_u0<=reg_1a8e23c7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0b346188_result_delayed_u0<=1'h0;
else reg_0b346188_result_delayed_u0<=reg_0b346188_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_11bf5a5d_u0<=1'h0;
else reg_11bf5a5d_u0<=reg_42f8ea27_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7b11510d_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_7b11510d_result_delayed_result_delayed_result_delayed_u0<=reg_7b11510d_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_16d553cc_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_16d553cc_result_delayed_result_delayed_result_delayed_u0<=reg_16d553cc_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4cf0ecf8_result_delayed_result_delayed_u0<=1'h0;
else reg_4cf0ecf8_result_delayed_result_delayed_u0<=reg_4cf0ecf8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_46180292_result_delayed_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_46180292_result_delayed_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_46180292_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1d5b7d72_result_delayed_result_delayed_u0<=1'h0;
else reg_1d5b7d72_result_delayed_result_delayed_u0<=reg_1d5b7d72_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2892d198_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_2892d198_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_2892d198_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_33d17fbe_result_delayed_result_delayed_u0<=1'h0;
else reg_33d17fbe_result_delayed_result_delayed_u0<=reg_33d17fbe_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7bbff74c_result_delayed_result_delayed_u0<=1'h0;
else reg_7bbff74c_result_delayed_result_delayed_u0<=reg_7bbff74c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4d591d1c_result_delayed_u0<=1'h0;
else reg_4d591d1c_result_delayed_u0<=reg_4d591d1c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u174<=1'h0;
else and_delayed_u174<=and_u2688_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2c350944_result_delayed_u0<=1'h0;
else reg_2c350944_result_delayed_u0<=reg_2c350944_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6ff6deb2_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_6ff6deb2_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_6ff6deb2_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2d137930_result_delayed_u0<=1'h0;
else reg_2d137930_result_delayed_u0<=reg_2d137930_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_42f8ea27_result_delayed_result_delayed_u0<=1'h0;
else reg_42f8ea27_result_delayed_result_delayed_u0<=reg_42f8ea27_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0a55fe82_result_delayed_result_delayed_u0<=1'h0;
else reg_0a55fe82_result_delayed_result_delayed_u0<=reg_0a55fe82_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_55043b64_result_delayed_u0<=1'h0;
else reg_55043b64_result_delayed_u0<=reg_55043b64_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_50915049_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_50915049_result_delayed_result_delayed_result_delayed_u0<=reg_50915049_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7c87d14d_result_delayed_u0<=1'h0;
else reg_7c87d14d_result_delayed_u0<=reg_7c87d14d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0c581759_u0<=1'h0;
else reg_0c581759_u0<=and_u2690_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3fcc3d8e_u0<=1'h0;
else reg_3fcc3d8e_u0<=reg_102f357e_result_delayed_result_delayed_u0;
end
assign or_u795_u0=reg_7b7cf4e5_u0|or_u793_u0;
assign or_u796_u0=and_u2690_u0|and_u2687_u0;
assign or_u797_u0=and_u2690_u0|and_u2687_u0;
assign or_u798_u0=and_u2690_u0|and_u2687_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_102f357e_u0<=1'h0;
else reg_102f357e_u0<=reg_0c581759_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7b7cf4e5_u0<=1'h0;
else reg_7b7cf4e5_u0<=reg_3fcc3d8e_result_delayed_u0;
end
assign and_u2689_u0=and_u2680_u0&and_u2691_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0c581759_result_delayed_u0<=1'h0;
else reg_0c581759_result_delayed_u0<=reg_0c581759_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3fcc3d8e_result_delayed_u0<=1'h0;
else reg_3fcc3d8e_result_delayed_u0<=reg_3fcc3d8e_u0;
end
assign and_u2690_u0=and_u2681_u0&and_u2691_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_102f357e_result_delayed_u0<=1'h0;
else reg_102f357e_result_delayed_u0<=reg_102f357e_u0;
end
assign or_u799_u0=and_u2690_u0|or_u794_u0;
assign mux_u271_u0=(and_u2690_u0)?1'h1:mux_u270;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0c581759_result_delayed_result_delayed_u0<=1'h0;
else reg_0c581759_result_delayed_result_delayed_u0<=reg_0c581759_result_delayed_u0;
end
assign or_u800_u0=and_u2690_u0|and_u2687_u0;
assign mux_u272_u0=(and_u2690_u0)?32'h8:32'h200;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_102f357e_result_delayed_result_delayed_u0<=1'h0;
else reg_102f357e_result_delayed_result_delayed_u0<=reg_102f357e_result_delayed_u0;
end
assign and_u2691_u0=and_u2678_u0&and_u2710_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6e7913b6_u0<=1'h0;
else reg_6e7913b6_u0<=and_u2692_u0;
end
assign or_u801_u0=or_u795_u0|reg_6e7913b6_u0;
assign and_u2692_u0=and_u2679_u0&and_u2710_u0;
assign equals_u142_a_signed={31'b0, port_7545a1a4_};
assign equals_u142_b_signed=32'h1;
assign equals_u142=equals_u142_a_signed==equals_u142_b_signed;
assign not_u470_u0=~equals_u142;
assign and_u2693_u0=and_u2710_u0&equals_u142;
assign and_u2694_u0=and_u2710_u0&not_u470_u0;
assign and_u2695_u0=and_u2709_u0&not_u471_u0;
assign and_u2696_u0=and_u2709_u0&port_05f8f754_;
assign not_u471_u0=~port_05f8f754_;
assign lessThan_u63_a_signed=port_1121f1ff_;
assign lessThan_u63_b_signed=port_70929f20_;
assign lessThan_u63=lessThan_u63_a_signed<lessThan_u63_b_signed;
assign and_u2697_u0=and_u2707_u0&lessThan_u63;
assign not_u472_u0=~lessThan_u63;
assign and_u2698_u0=and_u2707_u0&not_u472_u0;
assign not_u473_u0=~port_5286b1a6_;
assign and_u2699_u0=and_u2705_u0&not_u473_u0;
assign and_u2700_u0=and_u2705_u0&port_5286b1a6_;
assign add=port_1121f1ff_+32'h0;
assign and_u2701_u0=and_u2702_u0&port_1f63f705_;
assign simplePinWrite_u418=port_0a0e1767_;
assign simplePinWrite_u419=and_u2702_u0&{1{and_u2702_u0}};
assign simplePinWrite_u420=16'h1&{16{1'h1}};
assign add_u272=port_1121f1ff_+32'h1;
always @(posedge CLK)
begin
if (and_u2702_u0)
syncEnable_u434<=port_0a0e1767_;
end
always @(posedge CLK)
begin
if (and_u2705_u0)
syncEnable_u435_u0<=mux_u284_u0;
end
assign and_u2702_u0=and_u2700_u0&and_u2705_u0;
assign and_u2703_u0=and_u2699_u0&and_u2705_u0;
assign mux_u273_u0=(and_delayed_u175_u0)?syncEnable_u434:syncEnable_u435_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u175_u0<=1'h0;
else and_delayed_u175_u0<=and_u2702_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u176_u0<=1'h0;
else and_delayed_u176_u0<=and_u2703_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0f183598_u0<=1'h0;
else reg_0f183598_u0<=and_u2704_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4418b1bb_u0<=1'h0;
else reg_4418b1bb_u0<=and_u2705_u0;
end
assign mux_u274_u0=(reg_4418b1bb_u0)?syncEnable_u436_u0:32'h0;
always @(posedge CLK)
begin
if (and_u2707_u0)
syncEnable_u436_u0<=mux_u285_u0;
end
assign and_u2704_u0=and_u2698_u0&and_u2707_u0;
always @(posedge CLK)
begin
if (and_u2707_u0)
syncEnable_u437_u0<=mux_u284_u0;
end
assign mux_u275_u0=(reg_4418b1bb_u0)?mux_u273_u0:syncEnable_u437_u0;
assign and_u2705_u0=and_u2697_u0&and_u2707_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_532d6b49_u0<=1'h0;
else reg_532d6b49_u0<=and_u2707_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0b4f0828_u0<=1'h0;
else reg_0b4f0828_u0<=and_u2706_u0;
end
always @(posedge CLK)
begin
if (and_u2709_u0)
syncEnable_u438_u0<=mux_u285_u0;
end
assign mux_u276_u0=(reg_0b4f0828_u0)?syncEnable_u439_u0:mux_u275_u0;
always @(posedge CLK)
begin
if (and_u2709_u0)
syncEnable_u439_u0<=mux_u284_u0;
end
assign mux_u277_u0=(reg_0b4f0828_u0)?syncEnable_u438_u0:mux_u274_u0;
assign and_u2706_u0=and_u2695_u0&and_u2709_u0;
assign and_u2707_u0=and_u2696_u0&and_u2709_u0;
assign and_u2708_u0=and_u2694_u0&and_u2710_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_67514dd2_u0<=1'h0;
else reg_67514dd2_u0<=and_u2709_u0;
end
assign mux_u278_u0=(and_delayed_u177_u0)?syncEnable_u440_u0:mux_u277_u0;
assign mux_u279_u0=(and_delayed_u177_u0)?syncEnable_u441_u0:mux_u276_u0;
always @(posedge CLK)
begin
if (and_u2710_u0)
syncEnable_u440_u0<=mux_u285_u0;
end
assign and_u2709_u0=and_u2693_u0&and_u2710_u0;
always @(posedge CLK)
begin
if (and_u2710_u0)
syncEnable_u441_u0<=mux_u284_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u177_u0<=1'h0;
else and_delayed_u177_u0<=and_u2708_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
block_GO_delayed_u9<=1'h0;
else block_GO_delayed_u9<=and_u2710_u0;
end
assign mux_u280_u0=(or_u799_u0)?mux_u271_u0:1'h0;
assign or_u802_u0=or_u799_u0|and_u2704_u0;
assign latch_06dfa717_out=(block_GO_delayed_u9)?mux_u278_u0:latch_06dfa717_reg;
always @(posedge CLK)
begin
if (block_GO_delayed_u9)
latch_06dfa717_reg<=mux_u278_u0;
end
always @(posedge CLK)
begin
if (block_GO_delayed_u9)
latch_577ad7b1_reg<=mux_u279_u0;
end
assign latch_577ad7b1_out=(block_GO_delayed_u9)?mux_u279_u0:latch_577ad7b1_reg;
assign mux_u281_u0=(or_u800_u0)?{22'b0, mux_u272_u0[9], 5'b0, mux_u272_u0[3], 3'b0}:32'hffffffff;
assign or_u803_u0=or_u800_u0|and_u2704_u0;
assign or_u804_u0=or_u798_u0|and_u2704_u0;
assign mux_u282_u0=(or_u798_u0)?1'h1:1'h0;
assign or_u805_u0=or_u797_u0|and_u2702_u0;
assign mux_u283_u0=(or_u797_u0)?32'h0:add_u272;
assign and_u2710_u0=or_u806_u0&or_u806_u0;
always @(posedge CLK)
begin
if (or_u801_u0)
fbReg_temp_fsmOldState_resized_HH3_xy_5_u0<=latch_06dfa717_out;
end
assign mux_u284_u0=(loopControl_u6)?fbReg_Out1Portvalue_u2:16'h0;
always @(posedge CLK)
begin
if (reg_6f91e613_result_delayed_u0)
syncEnable_u442_u0<=RESET;
end
always @(posedge CLK)
begin
if (or_u801_u0)
fbReg_Out1Portvalue_u2<=latch_577ad7b1_out;
end
assign or_u806_u0=loopControl_u6|reg_6f91e613_result_delayed_u0;
assign mux_u285_u0=(loopControl_u6)?fbReg_temp_fsmOldState_resized_HH3_xy_5_u0:32'h0;
always @(posedge CLK or posedge syncEnable_u442_u0)
begin
if (syncEnable_u442_u0)
loopControl_u6<=1'h0;
else loopControl_u6<=or_u801_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6f91e613_u0<=1'h0;
else reg_6f91e613_u0<=GO;
end
assign mux_u286_u0=(GO)?32'h0:mux_u283_u0;
assign or_u807_u0=GO|or_u805_u0;
assign or_u808_u0=GO|or_u803_u0;
assign mux_u287_u0=(GO)?32'hffffffff:mux_u281_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6f91e613_result_delayed_u0<=1'h0;
else reg_6f91e613_result_delayed_u0<=reg_6f91e613_u0;
end
assign or_u809_u0=GO|or_u802_u0;
assign mux_u288_u0=(GO)?1'h0:mux_u280_u0;
assign or_u810_u0=GO|or_u804_u0;
assign mux_u289_u0=(GO)?1'h0:mux_u282_u0;
assign or_u811_u0=GO|or_u796_u0;
assign RESULT=or_u811_u0;
assign RESULT_u1604=32'h0;
assign RESULT_u1605=or_u809_u0;
assign RESULT_u1606=mux_u288_u0;
assign RESULT_u1607=or_u807_u0;
assign RESULT_u1608=mux_u286_u0;
assign RESULT_u1609=or_u808_u0;
assign RESULT_u1610=mux_u287_u0;
assign RESULT_u1611=or_u810_u0;
assign RESULT_u1612=mux_u289_u0;
assign RESULT_u1613=and_u2702_u0;
assign RESULT_u1614=add;
assign RESULT_u1615=3'h1;
assign RESULT_u1616=simplePinWrite_u419;
assign RESULT_u1617=simplePinWrite_u420;
assign RESULT_u1618=simplePinWrite_u417;
assign RESULT_u1619=simplePinWrite;
assign RESULT_u1620=simplePinWrite_u418;
assign RESULT_u1621=simplePinWrite_u416;
assign DONE=1'h0;
endmodule



module resized_HH3_xy_endianswapper_01d48b74_(endianswapper_01d48b74_in, endianswapper_01d48b74_out);
input	[31:0]	endianswapper_01d48b74_in;
output	[31:0]	endianswapper_01d48b74_out;
assign endianswapper_01d48b74_out=32'h0;
endmodule



module resized_HH3_xy_endianswapper_1a227e6d_(endianswapper_1a227e6d_in, endianswapper_1a227e6d_out);
input	[31:0]	endianswapper_1a227e6d_in;
output	[31:0]	endianswapper_1a227e6d_out;
assign endianswapper_1a227e6d_out=32'h0;
endmodule



module resized_HH3_xy_stateVar_fsmOldState_resized_HH3_xy(bus_265f821d_, bus_15b24ce3_, bus_4cadd642_, bus_11ea79c0_, bus_02dad7ef_);
input		bus_265f821d_;
input		bus_15b24ce3_;
input		bus_4cadd642_;
input	[31:0]	bus_11ea79c0_;
output	[31:0]	bus_02dad7ef_;
wire	[31:0]	endianswapper_01d48b74_out;
wire	[31:0]	endianswapper_1a227e6d_out;
resized_HH3_xy_endianswapper_01d48b74_ resized_HH3_xy_endianswapper_01d48b74__1(.endianswapper_01d48b74_in(32'h0), 
  .endianswapper_01d48b74_out(endianswapper_01d48b74_out));
assign bus_02dad7ef_=32'h0;
resized_HH3_xy_endianswapper_1a227e6d_ resized_HH3_xy_endianswapper_1a227e6d__1(.endianswapper_1a227e6d_in(32'h0), 
  .endianswapper_1a227e6d_out(endianswapper_1a227e6d_out));
endmodule



module resized_HH3_xy_endianswapper_1e4fe208_(endianswapper_1e4fe208_in, endianswapper_1e4fe208_out);
input	[31:0]	endianswapper_1e4fe208_in;
output	[31:0]	endianswapper_1e4fe208_out;
assign endianswapper_1e4fe208_out=endianswapper_1e4fe208_in;
endmodule



module resized_HH3_xy_endianswapper_3b262bed_(endianswapper_3b262bed_in, endianswapper_3b262bed_out);
input	[31:0]	endianswapper_3b262bed_in;
output	[31:0]	endianswapper_3b262bed_out;
assign endianswapper_3b262bed_out=endianswapper_3b262bed_in;
endmodule



module resized_HH3_xy_stateVar_Out1MaxTokenIndex(bus_24944e90_, bus_67a2773e_, bus_4329e6b2_, bus_31a05489_, bus_6ec88e4d_);
input		bus_24944e90_;
input		bus_67a2773e_;
input		bus_4329e6b2_;
input	[31:0]	bus_31a05489_;
output	[31:0]	bus_6ec88e4d_;
wire	[31:0]	endianswapper_1e4fe208_out;
reg	[31:0]	stateVar_Out1MaxTokenIndex_u2=32'h0;
wire	[31:0]	endianswapper_3b262bed_out;
resized_HH3_xy_endianswapper_1e4fe208_ resized_HH3_xy_endianswapper_1e4fe208__1(.endianswapper_1e4fe208_in(bus_31a05489_), 
  .endianswapper_1e4fe208_out(endianswapper_1e4fe208_out));
assign bus_6ec88e4d_=endianswapper_3b262bed_out;
always @(posedge bus_24944e90_ or posedge bus_67a2773e_)
begin
if (bus_67a2773e_)
stateVar_Out1MaxTokenIndex_u2<=32'h0;
else if (bus_4329e6b2_)
stateVar_Out1MaxTokenIndex_u2<=endianswapper_1e4fe208_out;
end
resized_HH3_xy_endianswapper_3b262bed_ resized_HH3_xy_endianswapper_3b262bed__1(.endianswapper_3b262bed_in(stateVar_Out1MaxTokenIndex_u2), 
  .endianswapper_3b262bed_out(endianswapper_3b262bed_out));
endmodule



module resized_HH3_xy_consumeRow(CLK, RESET, GO, port_36ed5a59_, port_55b6d605_, port_7a6b4a4c_, port_6b0ac5ca_, RESULT, RESULT_u1622, RESULT_u1623, RESULT_u1624, RESULT_u1625, RESULT_u1626, RESULT_u1627, RESULT_u1628, RESULT_u1629, RESULT_u1630, RESULT_u1631, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_36ed5a59_;
input		port_55b6d605_;
input		port_7a6b4a4c_;
input	[15:0]	port_6b0ac5ca_;
output		RESULT;
output	[15:0]	RESULT_u1622;
output		RESULT_u1623;
output	[31:0]	RESULT_u1624;
output	[15:0]	RESULT_u1625;
output	[2:0]	RESULT_u1626;
output		RESULT_u1627;
output	[31:0]	RESULT_u1628;
output	[15:0]	RESULT_u1629;
output	[2:0]	RESULT_u1630;
output		RESULT_u1631;
output		DONE;
wire		simplePinWrite;
wire		and_u2711_u0;
wire	[31:0]	add;
wire	[31:0]	add_u273;
wire		and_u2712_u0;
reg		reg_6459225d_u0=1'h0;
wire		or_u812_u0;
wire	[15:0]	add_u274;
reg	[15:0]	syncEnable_u443=16'h0;
wire		and_u2713_u0;
reg		and_delayed_u178=1'h0;
wire		lessThanEqualTo;
wire signed	[16:0]	lessThanEqualTo_a_signed;
wire signed	[16:0]	lessThanEqualTo_b_signed;
wire		and_u2714_u0;
wire		not_u474_u0;
wire		and_u2715_u0;
wire	[15:0]	mux_u290;
wire	[15:0]	latch_6301f4e8_out;
reg	[15:0]	latch_6301f4e8_reg=16'h0;
wire		or_u813_u0;
wire	[15:0]	add_u275;
wire		and_u2716_u0;
wire signed	[16:0]	lessThanEqualTo_u2_a_signed;
wire signed	[16:0]	lessThanEqualTo_u2_b_signed;
wire		lessThanEqualTo_u2;
wire		not_u475_u0;
wire		and_u2717_u0;
wire		and_u2718_u0;
wire	[15:0]	subtract;
wire	[31:0]	add_u276;
reg		reg_6e05f845_u0=1'h0;
wire		or_u814_u0;
wire		and_u2719_u0;
wire	[15:0]	add_u277;
reg	[15:0]	syncEnable_u444_u0=16'h0;
reg		reg_4ad5d3ee_u0=1'h0;
wire		and_u2720_u0;
reg	[15:0]	latch_1b9e3991_reg=16'h0;
wire	[15:0]	latch_1b9e3991_out;
wire	[15:0]	mux_u291_u0;
wire		or_u815_u0;
reg		reg_56a124c9_u0=1'h0;
reg	[15:0]	syncEnable_u445_u0=16'h0;
assign simplePinWrite=GO&{1{GO}};
assign and_u2711_u0=and_u2714_u0&or_u813_u0;
assign add={13'b0, port_36ed5a59_, 3'b0}+{mux_u290[15], mux_u290[15], mux_u290[15], mux_u290[15], mux_u290[15], mux_u290[15], mux_u290[15], mux_u290[15], mux_u290[15], mux_u290[15], mux_u290[15], mux_u290[15], mux_u290[15], mux_u290[15], mux_u290[15], mux_u290[15], mux_u290};
assign add_u273={add[20], add[20], add[20], add[20], add[20], add[20], add[20], add[20], add[20], add[20], add[20], add[20:0]}+32'h0;
assign and_u2712_u0=reg_6459225d_u0&port_55b6d605_;
always @(posedge CLK or posedge and_u2713_u0 or posedge or_u812_u0)
begin
if (or_u812_u0)
reg_6459225d_u0<=1'h0;
else if (and_u2713_u0)
reg_6459225d_u0<=1'h1;
else reg_6459225d_u0<=reg_6459225d_u0;
end
assign or_u812_u0=and_u2712_u0|RESET;
assign add_u274=mux_u290+16'h1;
always @(posedge CLK)
begin
if (and_u2713_u0)
syncEnable_u443<=add_u274;
end
assign and_u2713_u0=and_u2715_u0&or_u813_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u178<=1'h0;
else and_delayed_u178<=and_u2713_u0;
end
assign lessThanEqualTo_a_signed={mux_u290[15], mux_u290};
assign lessThanEqualTo_b_signed=17'h7;
assign lessThanEqualTo=lessThanEqualTo_a_signed<=lessThanEqualTo_b_signed;
assign and_u2714_u0=or_u813_u0&not_u474_u0;
assign not_u474_u0=~lessThanEqualTo;
assign and_u2715_u0=or_u813_u0&lessThanEqualTo;
assign mux_u290=(GO)?16'h0:syncEnable_u443;
assign latch_6301f4e8_out=(GO)?port_6b0ac5ca_:latch_6301f4e8_reg;
always @(posedge CLK)
begin
if (GO)
latch_6301f4e8_reg<=port_6b0ac5ca_;
end
assign or_u813_u0=GO|and_delayed_u178;
assign add_u275=port_36ed5a59_+16'h1;
assign and_u2716_u0=and_u2717_u0&or_u815_u0;
assign lessThanEqualTo_u2_a_signed={mux_u291_u0[15], mux_u291_u0};
assign lessThanEqualTo_u2_b_signed=17'h8;
assign lessThanEqualTo_u2=lessThanEqualTo_u2_a_signed<=lessThanEqualTo_u2_b_signed;
assign not_u475_u0=~lessThanEqualTo_u2;
assign and_u2717_u0=or_u815_u0&not_u475_u0;
assign and_u2718_u0=or_u815_u0&lessThanEqualTo_u2;
assign subtract=mux_u291_u0-16'h1;
assign add_u276={subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract}+32'h0;
always @(posedge CLK or posedge and_u2720_u0 or posedge or_u814_u0)
begin
if (or_u814_u0)
reg_6e05f845_u0<=1'h0;
else if (and_u2720_u0)
reg_6e05f845_u0<=1'h1;
else reg_6e05f845_u0<=reg_6e05f845_u0;
end
assign or_u814_u0=and_u2719_u0|RESET;
assign and_u2719_u0=reg_6e05f845_u0&port_7a6b4a4c_;
assign add_u277=mux_u291_u0+16'h1;
always @(posedge CLK)
begin
if (and_u2720_u0)
syncEnable_u444_u0<=add_u277;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4ad5d3ee_u0<=1'h0;
else reg_4ad5d3ee_u0<=and_u2720_u0;
end
assign and_u2720_u0=and_u2718_u0&or_u815_u0;
always @(posedge CLK)
begin
if (GO)
latch_1b9e3991_reg<=port_6b0ac5ca_;
end
assign latch_1b9e3991_out=(GO)?port_6b0ac5ca_:latch_1b9e3991_reg;
assign mux_u291_u0=(reg_4ad5d3ee_u0)?syncEnable_u444_u0:16'h1;
assign or_u815_u0=reg_4ad5d3ee_u0|GO;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_56a124c9_u0<=1'h0;
else reg_56a124c9_u0<=and_u2711_u0;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u445_u0<=add_u275;
end
assign RESULT=and_u2711_u0;
assign RESULT_u1622=syncEnable_u445_u0;
assign RESULT_u1623=and_u2713_u0;
assign RESULT_u1624=add_u273;
assign RESULT_u1625=latch_6301f4e8_out;
assign RESULT_u1626=3'h1;
assign RESULT_u1627=and_u2720_u0;
assign RESULT_u1628=add_u276;
assign RESULT_u1629=latch_1b9e3991_out;
assign RESULT_u1630=3'h1;
assign RESULT_u1631=simplePinWrite;
assign DONE=reg_56a124c9_u0;
endmodule



module resized_HH3_xy_structuralmemory_068f5fb6_(CLK_u15, bus_13f3e3d1_, bus_750d9e9a_, bus_0cd70fa4_, bus_30fff37e_, bus_2ba929a7_, bus_6b58816e_, bus_035cdb42_, bus_1dbe1e5d_);
input		CLK_u15;
input		bus_13f3e3d1_;
input	[31:0]	bus_750d9e9a_;
input	[2:0]	bus_0cd70fa4_;
input		bus_30fff37e_;
input		bus_2ba929a7_;
input	[15:0]	bus_6b58816e_;
output	[15:0]	bus_035cdb42_;
output		bus_1dbe1e5d_;
wire		and_236dfa8f_u0;
wire		not_0537599c_u0;
reg		logicalMem_2a36bc10_we_delay0_u0=1'h0;
wire	[15:0]	bus_64d59103_;
wire		or_279802cd_u0;
wire		or_58a1523b_u0;
assign and_236dfa8f_u0=bus_30fff37e_&not_0537599c_u0;
assign not_0537599c_u0=~bus_2ba929a7_;
always @(posedge CLK_u15 or posedge bus_13f3e3d1_)
begin
if (bus_13f3e3d1_)
logicalMem_2a36bc10_we_delay0_u0<=1'h0;
else logicalMem_2a36bc10_we_delay0_u0<=bus_2ba929a7_;
end
assign bus_035cdb42_=bus_64d59103_;
assign bus_1dbe1e5d_=or_279802cd_u0;
resized_HH3_xy_forge_memory_512x16_28 resized_HH3_xy_forge_memory_512x16_28_instance1(.CLK(CLK_u15), 
  .EN(or_58a1523b_u0), .WE(bus_2ba929a7_), .ADDR(bus_750d9e9a_), .DIN(bus_6b58816e_), 
  .DOUT(bus_64d59103_), .DONE());
assign or_279802cd_u0=and_236dfa8f_u0|logicalMem_2a36bc10_we_delay0_u0;
assign or_58a1523b_u0=bus_30fff37e_|bus_2ba929a7_;
endmodule


