// __  ___ __ ___  _ __   ___  ___ 
// \ \/ / '__/ _ \| '_ \ / _ \/ __|
//  >  <| | | (_) | | | | (_) \__ \
// /_/\_\_|  \___/|_| |_|\___/|___/
// 
// Xronos synthesizer version
// Run date: Thu 2 Nov 2017 13:56:10 +0000
// 

module LL1_H_iunzipFilter2D(In1_DATA, In1_SEND, Out2_DATA, Out2_COUNT, Out1_ACK, In1_ACK, Out2_ACK, Out1_RDY, Out1_COUNT, Out2_RDY, CLK, Out2_SEND, Out1_SEND, Out1_DATA, RESET, In1_COUNT);
wire		topRow_go;
input	[15:0]	In1_DATA;
wire		midNoConsume1_go;
input		In1_SEND;
wire		mid2_go;
wire		bottomLeftNoConsume1_done;
wire		bottomRightNoConsume2_done;
output	[15:0]	Out2_DATA;
wire		bottomRowNoConsume1_go;
wire		midLeftNoConsume2_done;
wire		bottomLeftNoConsume1_go;
wire		midLeft1_done;
wire		midNoConsume2_done;
wire		bottomRowNoConsume2_go;
wire		topRight_done;
wire		populateBuffer_go;
wire		midRight2_done;
output	[15:0]	Out2_COUNT;
wire		populateBuffer_done;
wire		bottomRightNoConsume1_go;
input		Out1_ACK;
output		In1_ACK;
wire		midLeft1_go;
wire		bottomRowNoConsume1_done;
wire		topRight_go;
wire		midLeftNoConsume2_go;
wire		bottomRightNoConsume2_go;
wire		midLeft2_done;
input		Out2_ACK;
wire		donePopulateBuffer_done;
input		Out1_RDY;
wire		topLeft_go;
wire		mid1_done;
wire		bottomLeftNoConsume2_done;
wire		bottomRightNoConsume1_done;
wire		midRightNoConsume1_go;
output	[15:0]	Out1_COUNT;
wire		midLeftNoConsume1_go;
input		Out2_RDY;
wire		midRight1_go;
wire		donePopulateBuffer_go;
wire		midNoConsume2_go;
wire		midRightNoConsume2_go;
input		CLK;
wire		topLeft_done;
wire		mid2_done;
wire		mid1_go;
wire		midNoConsume1_done;
wire		midRight2_go;
output		Out2_SEND;
wire		bottomRowNoConsume2_done;
output		Out1_SEND;
wire		midLeft2_go;
wire		midRightNoConsume1_done;
output	[15:0]	Out1_DATA;
input		RESET;
wire		topRow_done;
input	[15:0]	In1_COUNT;
wire		midLeftNoConsume1_done;
wire		midRight1_done;
wire		bottomLeftNoConsume2_go;
wire		midRightNoConsume2_done;
wire		LL1_H_iunzipFilter2D_midLeftNoConsume1_instance_DONE;
wire	[15:0]	midLeftNoConsume1_u8;
wire	[15:0]	midLeftNoConsume1_u6;
wire	[15:0]	midLeftNoConsume1_u0;
wire		midLeftNoConsume1_u7;
wire	[31:0]	midLeftNoConsume1_u4;
wire		midLeftNoConsume1_u3;
wire	[15:0]	midLeftNoConsume1_u2;
wire	[2:0]	midLeftNoConsume1_u5;
wire		midLeftNoConsume1;
wire		midLeftNoConsume1_u1;
wire		bus_7c830cee_;
wire		bottomRowNoConsume1;
wire	[15:0]	bottomRowNoConsume1_u0;
wire	[31:0]	bottomRowNoConsume1_u4;
wire		LL1_H_iunzipFilter2D_bottomRowNoConsume1_instance_DONE;
wire		bottomRowNoConsume1_u1;
wire	[15:0]	bottomRowNoConsume1_u2;
wire		bottomRowNoConsume1_u3;
wire	[2:0]	bottomRowNoConsume1_u5;
wire	[15:0]	bottomRowNoConsume1_u6;
wire		bottomRowNoConsume1_u7;
wire	[15:0]	bottomRowNoConsume1_u8;
wire		bus_47e0da85_;
wire		bus_279a0f63_;
wire		midRightNoConsume2_u3;
wire		midRightNoConsume2;
wire		midRightNoConsume2_u1;
wire		midRightNoConsume2_u4;
wire	[2:0]	midRightNoConsume2_u7;
wire	[15:0]	midRightNoConsume2_u8;
wire		midRightNoConsume2_u5;
wire	[31:0]	midRightNoConsume2_u6;
wire	[15:0]	midRightNoConsume2_u2;
wire	[15:0]	midRightNoConsume2_u0;
wire		midRightNoConsume2_u10;
wire	[15:0]	midRightNoConsume2_u9;
wire		LL1_H_iunzipFilter2D_midRightNoConsume2_instance_DONE;
wire		bottomLeftNoConsume1_u7;
wire	[15:0]	bottomLeftNoConsume1_u8;
wire	[2:0]	bottomLeftNoConsume1_u5;
wire		LL1_H_iunzipFilter2D_bottomLeftNoConsume1_instance_DONE;
wire	[15:0]	bottomLeftNoConsume1_u2;
wire	[15:0]	bottomLeftNoConsume1_u6;
wire		bottomLeftNoConsume1;
wire	[15:0]	bottomLeftNoConsume1_u0;
wire		bottomLeftNoConsume1_u3;
wire		bottomLeftNoConsume1_u1;
wire	[31:0]	bottomLeftNoConsume1_u4;
wire		bus_0f1f6bab_;
wire	[15:0]	mid1_u15;
wire	[2:0]	mid1_u11;
wire		mid1_u12;
wire	[15:0]	mid1_u2;
wire		mid1_u9;
wire		mid1_u3;
wire	[15:0]	mid1_u4;
wire	[2:0]	mid1_u8;
wire		mid1_u5;
wire	[31:0]	mid1_u6;
wire	[31:0]	mid1_u10;
wire		mid1;
wire	[31:0]	mid1_u0;
wire		mid1_u1;
wire	[15:0]	mid1_u7;
wire		LL1_H_iunzipFilter2D_mid1_instance_DONE;
wire		mid1_u14;
wire	[15:0]	mid1_u13;
wire		midLeftNoConsume2_u7;
wire	[15:0]	midLeftNoConsume2_u6;
wire		LL1_H_iunzipFilter2D_midLeftNoConsume2_instance_DONE;
wire		midLeftNoConsume2_u3;
wire		midLeftNoConsume2;
wire	[15:0]	midLeftNoConsume2_u0;
wire	[15:0]	midLeftNoConsume2_u2;
wire	[31:0]	midLeftNoConsume2_u4;
wire	[15:0]	midLeftNoConsume2_u8;
wire	[2:0]	midLeftNoConsume2_u5;
wire		midLeftNoConsume2_u1;
wire		bus_1564633b_;
wire	[15:0]	bus_5ad36c45_;
wire		bus_7a837774_;
wire		bus_15ecd674_;
wire		or_396b3042_u0;
wire	[15:0]	bus_7d411a66_;
wire		bus_3fffd7cb_;
wire	[31:0]	bus_2da7af10_;
wire		bus_624df4b1_;
wire	[2:0]	bus_77051f23_;
wire		bus_3681a366_;
wire		LL1_H_iunzipFilter2D_midLeft1_instance_DONE;
wire		midLeft1_u9;
wire		midLeft1;
wire	[15:0]	midLeft1_u4;
wire	[15:0]	midLeft1_u15;
wire	[2:0]	midLeft1_u11;
wire		midLeft1_u12;
wire	[15:0]	midLeft1_u7;
wire	[31:0]	midLeft1_u10;
wire	[2:0]	midLeft1_u8;
wire	[31:0]	midLeft1_u2;
wire		midLeft1_u3;
wire		midLeft1_u5;
wire	[31:0]	midLeft1_u6;
wire		midLeft1_u14;
wire	[15:0]	midLeft1_u0;
wire		midLeft1_u1;
wire	[15:0]	midLeft1_u13;
wire		bus_0379aee9_;
wire		bus_73d09570_;
wire		bus_4ae3b466_;
wire		or_0823cb19_u0;
wire		bus_52c37c26_;
wire		bus_46448f94_;
wire		bus_12ce21da_;
wire		bus_5d6bea1c_;
wire		bus_4f3a32a9_;
wire		donePopulateBuffer;
wire	[15:0]	donePopulateBuffer_u0;
wire		LL1_H_iunzipFilter2D_donePopulateBuffer_instance_DONE;
wire	[2:0]	bus_60d84d20_;
wire	[15:0]	or_76a627f2_u0;
wire		bus_4ca9c49f_;
wire	[15:0]	bottomRightNoConsume1_u12;
wire	[15:0]	bottomRightNoConsume1_u4;
wire		bottomRightNoConsume1_u3;
wire		bottomRightNoConsume1_u1;
wire	[2:0]	bottomRightNoConsume1_u11;
wire		bottomRightNoConsume1;
wire		LL1_H_iunzipFilter2D_bottomRightNoConsume1_instance_DONE;
wire		bottomRightNoConsume1_u9;
wire	[15:0]	bottomRightNoConsume1_u14;
wire		bottomRightNoConsume1_u13;
wire		bottomRightNoConsume1_u7;
wire		bottomRightNoConsume1_u5;
wire	[31:0]	bottomRightNoConsume1_u10;
wire		bottomRightNoConsume1_u8;
wire	[15:0]	bottomRightNoConsume1_u2;
wire	[15:0]	bottomRightNoConsume1_u0;
wire	[31:0]	bottomRightNoConsume1_u6;
wire		bus_15ebb497_;
wire	[15:0]	bottomLeftNoConsume2_u6;
wire		bottomLeftNoConsume2_u7;
wire		LL1_H_iunzipFilter2D_bottomLeftNoConsume2_instance_DONE;
wire	[2:0]	bottomLeftNoConsume2_u5;
wire		bottomLeftNoConsume2_u3;
wire		bottomLeftNoConsume2;
wire		bottomLeftNoConsume2_u1;
wire	[15:0]	bottomLeftNoConsume2_u8;
wire	[15:0]	bottomLeftNoConsume2_u0;
wire	[15:0]	bottomLeftNoConsume2_u2;
wire	[31:0]	bottomLeftNoConsume2_u4;
wire		topLeft;
wire	[31:0]	topLeft_u6;
wire	[15:0]	topLeft_u0;
wire		topLeft_u3;
wire		topLeft_u5;
wire		topLeft_u12;
wire		topLeft_u14;
wire	[31:0]	topLeft_u9;
wire	[2:0]	topLeft_u11;
wire	[2:0]	topLeft_u7;
wire	[15:0]	topLeft_u4;
wire	[15:0]	topLeft_u10;
wire	[15:0]	topLeft_u13;
wire	[31:0]	topLeft_u2;
wire	[15:0]	topLeft_u15;
wire		LL1_H_iunzipFilter2D_topLeft_instance_DONE;
wire		topLeft_u1;
wire		topLeft_u8;
wire		topRight_u18;
wire	[15:0]	topRight_u19;
wire	[15:0]	topRight_u6;
wire	[2:0]	topRight_u11;
wire	[15:0]	topRight_u17;
wire	[31:0]	topRight_u13;
wire		topRight_u1;
wire	[2:0]	topRight_u15;
wire		topRight;
wire	[31:0]	topRight_u0;
wire		topRight_u3;
wire		topRight_u5;
wire	[15:0]	topRight_u2;
wire	[15:0]	topRight_u14;
wire		topRight_u16;
wire	[15:0]	topRight_u4;
wire		topRight_u12;
wire		topRight_u7;
wire		LL1_H_iunzipFilter2D_topRight_instance_DONE;
wire		topRight_u9;
wire		topRight_u8;
wire	[31:0]	topRight_u10;
wire	[15:0]	bus_25361c61_;
wire	[15:0]	bus_6dd7c8fd_;
wire		bus_7faecdeb_;
wire		bus_02cec1f3_;
wire	[15:0]	midNoConsume1_u8;
wire	[15:0]	midNoConsume1_u0;
wire	[15:0]	midNoConsume1_u2;
wire		midNoConsume1_u3;
wire	[31:0]	midNoConsume1_u4;
wire		midNoConsume1_u7;
wire		midNoConsume1;
wire	[15:0]	midNoConsume1_u6;
wire	[2:0]	midNoConsume1_u5;
wire		midNoConsume1_u1;
wire		LL1_H_iunzipFilter2D_midNoConsume1_instance_DONE;
wire	[15:0]	midNoConsume2_u6;
wire		midNoConsume2_u3;
wire		midNoConsume2_u8;
wire		LL1_H_iunzipFilter2D_midNoConsume2_instance_DONE;
wire	[15:0]	midNoConsume2_u2;
wire	[31:0]	midNoConsume2_u4;
wire		midNoConsume2_u1;
wire	[15:0]	midNoConsume2_u0;
wire	[15:0]	midNoConsume2_u7;
wire		midNoConsume2;
wire	[2:0]	midNoConsume2_u5;
wire		bus_1f82e86b_;
wire	[15:0]	or_0315d09f_u0;
wire		bus_6f5c9bce_;
wire		bus_386c7386_;
wire	[15:0]	bus_42424c02_;
wire	[15:0]	bus_35bb43c2_;
wire	[15:0]	bus_02c8854d_;
wire	[15:0]	bus_6308ab98_;
wire	[15:0]	bus_5a1ddee7_;
wire	[15:0]	bus_1807f3cd_;
wire	[31:0]	bus_1446f926_;
wire	[15:0]	bus_27d78a2b_;
wire		bus_1f5c5926_;
wire	[15:0]	bus_2f7aa6e4_;
wire	[15:0]	bus_4b3e6981_;
wire	[15:0]	bus_5a5f2961_;
wire		bus_31710b5f_;
wire	[15:0]	bus_29c7540a_;
wire		bus_299c5c34_;
wire	[15:0]	bus_7b6d2db0_;
wire		bus_7e378a50_;
wire	[15:0]	bus_2c656446_;
wire		bus_75734968_;
wire		bus_78fb14d7_;
wire	[15:0]	bus_623e353f_;
wire		bus_782a49ae_;
wire		bus_0ad99597_;
wire		bus_1df60b90_;
wire	[2:0]	bus_4ad1a98a_;
wire		bus_018f435a_;
wire		bus_78addd53_;
wire		bus_05553665_;
wire	[15:0]	bus_03a2926d_;
wire	[15:0]	bus_12066278_;
wire		bus_3b77c854_;
wire	[15:0]	bus_5727ff78_;
wire	[15:0]	bus_167da5bd_;
wire		bus_57083dd4_;
wire		bus_0fd98caa_;
wire		bus_24ac86a8_;
wire		bus_5122026c_;
wire		bus_15fa8b31_;
wire	[15:0]	bus_13a61289_;
wire		bus_7b461753_;
wire	[15:0]	bus_7cd6911c_;
wire		bus_2781fc25_;
wire		bus_6341aa95_;
wire		bus_295fc32e_;
wire	[15:0]	bus_75b6e6aa_;
wire	[15:0]	bus_52935bd9_;
wire		bus_47b6d4cf_;
wire		topRow_u16;
wire		topRow_u14;
wire	[15:0]	topRow_u15;
wire	[15:0]	topRow_u6;
wire	[15:0]	topRow_u17;
wire	[31:0]	topRow_u8;
wire	[15:0]	topRow_u4;
wire	[2:0]	topRow_u13;
wire		topRow;
wire		topRow_u3;
wire		LL1_H_iunzipFilter2D_topRow_instance_DONE;
wire		topRow_u10;
wire	[31:0]	topRow_u11;
wire		topRow_u5;
wire	[15:0]	topRow_u2;
wire		topRow_u1;
wire	[31:0]	topRow_u0;
wire	[2:0]	topRow_u9;
wire		topRow_u7;
wire	[15:0]	topRow_u12;
wire	[15:0]	bus_2a7d4abb_;
wire	[2:0]	midRight2_u11;
wire	[15:0]	midRight2_u19;
wire		midRight2_u7;
wire		midRight2_u3;
wire	[15:0]	midRight2_u6;
wire		midRight2_u8;
wire		midRight2_u5;
wire		midRight2_u12;
wire	[15:0]	midRight2_u14;
wire	[2:0]	midRight2_u15;
wire		midRight2_u1;
wire	[31:0]	midRight2_u2;
wire	[31:0]	midRight2_u13;
wire		midRight2_u16;
wire		midRight2_u18;
wire		midRight2;
wire		midRight2_u9;
wire	[15:0]	midRight2_u4;
wire	[31:0]	midRight2_u10;
wire	[15:0]	midRight2_u17;
wire		LL1_H_iunzipFilter2D_midRight2_instance_DONE;
wire	[15:0]	midRight2_u0;
wire	[15:0]	or_31aa5212_u0;
wire		bus_23506230_;
wire	[15:0]	or_71cb5f0a_u0;
wire	[15:0]	bus_4cb9b263_;
wire		bus_67323e98_;
wire		bus_6f12b7f2_;
wire		bottomRightNoConsume2_u3;
wire	[31:0]	bottomRightNoConsume2_u10;
wire	[15:0]	bottomRightNoConsume2_u4;
wire		bottomRightNoConsume2_u5;
wire	[15:0]	bottomRightNoConsume2_u0;
wire		bottomRightNoConsume2_u1;
wire		bottomRightNoConsume2;
wire		bottomRightNoConsume2_u9;
wire	[15:0]	bottomRightNoConsume2_u12;
wire	[15:0]	bottomRightNoConsume2_u14;
wire		bottomRightNoConsume2_u13;
wire		LL1_H_iunzipFilter2D_bottomRightNoConsume2_instance_DONE;
wire		bottomRightNoConsume2_u7;
wire	[15:0]	bottomRightNoConsume2_u2;
wire	[31:0]	bottomRightNoConsume2_u6;
wire	[2:0]	bottomRightNoConsume2_u11;
wire		bottomRightNoConsume2_u8;
wire		mid2_u12;
wire	[15:0]	mid2_u2;
wire	[2:0]	mid2_u8;
wire		mid2_u9;
wire	[15:0]	mid2_u14;
wire	[31:0]	mid2_u10;
wire		mid2_u5;
wire		LL1_H_iunzipFilter2D_mid2_instance_DONE;
wire		mid2_u15;
wire	[31:0]	mid2_u6;
wire	[15:0]	mid2_u13;
wire	[31:0]	mid2_u0;
wire	[15:0]	mid2_u4;
wire	[2:0]	mid2_u11;
wire		mid2;
wire		mid2_u3;
wire	[15:0]	mid2_u7;
wire		mid2_u1;
wire	[15:0]	bottomRowNoConsume2_u0;
wire		bottomRowNoConsume2_u1;
wire	[15:0]	bottomRowNoConsume2_u6;
wire		LL1_H_iunzipFilter2D_bottomRowNoConsume2_instance_DONE;
wire	[15:0]	bottomRowNoConsume2_u2;
wire	[2:0]	bottomRowNoConsume2_u5;
wire		bottomRowNoConsume2_u3;
wire	[31:0]	bottomRowNoConsume2_u4;
wire		bottomRowNoConsume2;
wire		bottomRowNoConsume2_u8;
wire	[15:0]	bottomRowNoConsume2_u7;
wire		bus_184376b1_;
wire		or_4b5f8e83_u0;
wire		bus_3fb35a7b_;
wire	[15:0]	midLeft2_u4;
wire		midLeft2_u5;
wire		midLeft2_u1;
wire		midLeft2;
wire	[15:0]	midLeft2_u7;
wire	[2:0]	midLeft2_u11;
wire		midLeft2_u9;
wire		midLeft2_u3;
wire		LL1_H_iunzipFilter2D_midLeft2_instance_DONE;
wire		midLeft2_u14;
wire		midLeft2_u12;
wire	[15:0]	midLeft2_u15;
wire	[31:0]	midLeft2_u6;
wire	[2:0]	midLeft2_u8;
wire	[15:0]	midLeft2_u0;
wire	[31:0]	midLeft2_u10;
wire	[15:0]	midLeft2_u13;
wire	[31:0]	midLeft2_u2;
wire	[31:0]	bus_69808cf7_;
wire	[15:0]	bus_70eb3e5c_;
wire	[31:0]	populateBuffer_u4;
wire	[15:0]	populateBuffer_u5;
wire		populateBuffer_u1;
wire		LL1_H_iunzipFilter2D_populateBuffer_instance_DONE;
wire	[31:0]	populateBuffer_u2;
wire		populateBuffer_u7;
wire		populateBuffer;
wire		populateBuffer_u3;
wire	[15:0]	populateBuffer_u0;
wire	[2:0]	populateBuffer_u6;
wire		scheduler_u31;
wire		scheduler_u21;
wire		scheduler_u29;
wire		scheduler_u36;
wire		scheduler_u41;
wire		scheduler_u26;
wire		scheduler_u32;
wire		scheduler_u19;
wire		scheduler_u40;
wire		scheduler_u23;
wire		scheduler_u25;
wire		scheduler_u39;
wire		scheduler_u38;
wire		scheduler_u20;
wire		scheduler_u27;
wire		scheduler_u37;
wire		scheduler_u28;
wire		scheduler_u22;
wire		scheduler_u33;
wire		scheduler;
wire		scheduler_u24;
wire	[2:0]	scheduler_u18;
wire		scheduler_u34;
wire		LL1_H_iunzipFilter2D_scheduler_instance_DONE;
wire		scheduler_u30;
wire		scheduler_u35;
wire	[2:0]	midRightNoConsume1_u7;
wire	[15:0]	midRightNoConsume1_u10;
wire	[15:0]	midRightNoConsume1_u0;
wire	[15:0]	midRightNoConsume1_u8;
wire		midRightNoConsume1_u9;
wire		midRightNoConsume1_u4;
wire		midRightNoConsume1_u3;
wire		midRightNoConsume1;
wire	[31:0]	midRightNoConsume1_u6;
wire		midRightNoConsume1_u1;
wire		LL1_H_iunzipFilter2D_midRightNoConsume1_instance_DONE;
wire		midRightNoConsume1_u5;
wire	[15:0]	midRightNoConsume1_u2;
wire		bus_22299860_;
wire	[15:0]	midRight1_u11;
wire		midRight1_u13;
wire	[2:0]	midRight1_u12;
wire		midRight1_u7;
wire	[15:0]	midRight1_u19;
wire		midRight1_u3;
wire	[31:0]	midRight1_u10;
wire	[15:0]	midRight1_u17;
wire		midRight1_u8;
wire	[31:0]	midRight1_u2;
wire		midRight1_u5;
wire		midRight1_u9;
wire		LL1_H_iunzipFilter2D_midRight1_instance_DONE;
wire	[15:0]	midRight1_u4;
wire		midRight1_u18;
wire	[2:0]	midRight1_u15;
wire		midRight1;
wire	[15:0]	midRight1_u0;
wire	[15:0]	midRight1_u6;
wire	[31:0]	midRight1_u14;
wire		midRight1_u1;
wire		midRight1_u16;
assign topRow_go=scheduler_u22;
assign midNoConsume1_go=scheduler_u24;
assign mid2_go=scheduler_u30;
assign bottomLeftNoConsume1_done=bus_7a837774_;
assign bottomRightNoConsume2_done=bus_3fb35a7b_;
assign Out2_DATA=or_0315d09f_u0;
assign bottomRowNoConsume1_go=scheduler_u20;
assign midLeftNoConsume2_done=bus_0379aee9_;
assign bottomLeftNoConsume1_go=scheduler_u25;
assign midLeft1_done=bus_67323e98_;
assign midNoConsume2_done=bus_1f82e86b_;
assign bottomRowNoConsume2_go=scheduler_u31;
assign topRight_done=bus_52c37c26_;
assign populateBuffer_go=scheduler_u36;
assign midRight2_done=bus_22299860_;
assign Out2_COUNT=or_76a627f2_u0;
assign populateBuffer_done=bus_47e0da85_;
assign bottomRightNoConsume1_go=scheduler_u34;
assign In1_ACK=or_396b3042_u0;
assign midLeft1_go=scheduler_u19;
assign bottomRowNoConsume1_done=bus_279a0f63_;
assign topRight_go=scheduler_u26;
assign midLeftNoConsume2_go=scheduler_u27;
assign bottomRightNoConsume2_go=scheduler_u29;
assign midLeft2_done=bus_6f12b7f2_;
assign donePopulateBuffer_done=bus_46448f94_;
assign topLeft_go=scheduler_u40;
assign mid1_done=bus_5d6bea1c_;
assign bottomLeftNoConsume2_done=bus_4ca9c49f_;
assign bottomRightNoConsume1_done=bus_0f1f6bab_;
assign midRightNoConsume1_go=scheduler_u33;
assign Out1_COUNT=or_71cb5f0a_u0;
assign midLeftNoConsume1_go=scheduler_u37;
assign midRight1_go=scheduler_u39;
assign donePopulateBuffer_go=scheduler_u41;
assign midNoConsume2_go=scheduler_u21;
assign midRightNoConsume2_go=scheduler_u23;
assign topLeft_done=bus_6f5c9bce_;
assign mid2_done=bus_4f3a32a9_;
assign mid1_go=scheduler_u32;
assign midNoConsume1_done=bus_386c7386_;
assign midRight2_go=scheduler_u38;
assign Out2_SEND=or_0823cb19_u0;
assign bottomRowNoConsume2_done=bus_1564633b_;
assign Out1_SEND=or_4b5f8e83_u0;
assign midLeft2_go=scheduler_u35;
assign midRightNoConsume1_done=bus_15ecd674_;
assign Out1_DATA=or_31aa5212_u0;
assign topRow_done=bus_7c830cee_;
assign midLeftNoConsume1_done=bus_73d09570_;
assign midRight1_done=bus_184376b1_;
assign bottomLeftNoConsume2_go=scheduler_u28;
assign midRightNoConsume2_done=bus_12ce21da_;
LL1_H_iunzipFilter2D_midLeftNoConsume1 LL1_H_iunzipFilter2D_midLeftNoConsume1_instance(.CLK(CLK), 
  .RESET(bus_23506230_), .GO(midLeftNoConsume1_go), .port_24c1e388_(16'h0), .port_3d7d2b97_(bus_5ad36c45_), 
  .port_4f846b64_(bus_31710b5f_), .port_325dd0f8_(bus_12066278_), .DONE(LL1_H_iunzipFilter2D_midLeftNoConsume1_instance_DONE), 
  .RESULT(midLeftNoConsume1), .RESULT_u60(midLeftNoConsume1_u0), .RESULT_u61(midLeftNoConsume1_u1), 
  .RESULT_u62(midLeftNoConsume1_u2), .RESULT_u63(midLeftNoConsume1_u3), .RESULT_u64(midLeftNoConsume1_u4), 
  .RESULT_u65(midLeftNoConsume1_u5), .RESULT_u66(midLeftNoConsume1_u6), .RESULT_u67(midLeftNoConsume1_u7), 
  .RESULT_u68(midLeftNoConsume1_u8));
assign bus_7c830cee_=LL1_H_iunzipFilter2D_topRow_instance_DONE&{1{LL1_H_iunzipFilter2D_topRow_instance_DONE}};
LL1_H_iunzipFilter2D_bottomRowNoConsume1 LL1_H_iunzipFilter2D_bottomRowNoConsume1_instance(.CLK(CLK), 
  .RESET(bus_23506230_), .GO(bottomRowNoConsume1_go), .port_72ef45b3_(bus_5ad36c45_), 
  .port_6163a4df_(bus_75734968_), .port_1df2cf41_(bus_4b3e6981_), .DONE(LL1_H_iunzipFilter2D_bottomRowNoConsume1_instance_DONE), 
  .RESULT(bottomRowNoConsume1), .RESULT_u69(bottomRowNoConsume1_u0), .RESULT_u70(bottomRowNoConsume1_u1), 
  .RESULT_u71(bottomRowNoConsume1_u2), .RESULT_u72(bottomRowNoConsume1_u3), .RESULT_u73(bottomRowNoConsume1_u4), 
  .RESULT_u74(bottomRowNoConsume1_u5), .RESULT_u75(bottomRowNoConsume1_u6), .RESULT_u76(bottomRowNoConsume1_u7), 
  .RESULT_u77(bottomRowNoConsume1_u8));
assign bus_47e0da85_=LL1_H_iunzipFilter2D_populateBuffer_instance_DONE&{1{LL1_H_iunzipFilter2D_populateBuffer_instance_DONE}};
assign bus_279a0f63_=LL1_H_iunzipFilter2D_bottomRowNoConsume1_instance_DONE&{1{LL1_H_iunzipFilter2D_bottomRowNoConsume1_instance_DONE}};
LL1_H_iunzipFilter2D_midRightNoConsume2 LL1_H_iunzipFilter2D_midRightNoConsume2_instance(.CLK(CLK), 
  .RESET(bus_23506230_), .GO(midRightNoConsume2_go), .port_461847e8_(bus_4cb9b263_), 
  .port_24a7300a_(bus_15ebb497_), .port_03e1c37e_(bus_15fa8b31_), .port_0d8191ee_(bus_2c656446_), 
  .DONE(LL1_H_iunzipFilter2D_midRightNoConsume2_instance_DONE), .RESULT(midRightNoConsume2), 
  .RESULT_u78(midRightNoConsume2_u0), .RESULT_u79(midRightNoConsume2_u1), .RESULT_u80(midRightNoConsume2_u2), 
  .RESULT_u81(midRightNoConsume2_u3), .RESULT_u82(midRightNoConsume2_u4), .RESULT_u83(midRightNoConsume2_u5), 
  .RESULT_u84(midRightNoConsume2_u6), .RESULT_u85(midRightNoConsume2_u7), .RESULT_u86(midRightNoConsume2_u8), 
  .RESULT_u87(midRightNoConsume2_u9), .RESULT_u88(midRightNoConsume2_u10));
LL1_H_iunzipFilter2D_bottomLeftNoConsume1 LL1_H_iunzipFilter2D_bottomLeftNoConsume1_instance(.CLK(CLK), 
  .RESET(bus_23506230_), .GO(bottomLeftNoConsume1_go), .port_47f3deda_(16'h0), 
  .port_01459c00_(bus_5ad36c45_), .port_4b02a40f_(bus_24ac86a8_), .port_5e56587d_(bus_29c7540a_), 
  .DONE(LL1_H_iunzipFilter2D_bottomLeftNoConsume1_instance_DONE), .RESULT(bottomLeftNoConsume1), 
  .RESULT_u89(bottomLeftNoConsume1_u0), .RESULT_u90(bottomLeftNoConsume1_u1), 
  .RESULT_u91(bottomLeftNoConsume1_u2), .RESULT_u92(bottomLeftNoConsume1_u3), 
  .RESULT_u93(bottomLeftNoConsume1_u4), .RESULT_u94(bottomLeftNoConsume1_u5), 
  .RESULT_u95(bottomLeftNoConsume1_u6), .RESULT_u96(bottomLeftNoConsume1_u7), 
  .RESULT_u97(bottomLeftNoConsume1_u8));
assign bus_0f1f6bab_=LL1_H_iunzipFilter2D_bottomRightNoConsume1_instance_DONE&{1{LL1_H_iunzipFilter2D_bottomRightNoConsume1_instance_DONE}};
LL1_H_iunzipFilter2D_mid1 LL1_H_iunzipFilter2D_mid1_instance(.CLK(CLK), .RESET(bus_23506230_), 
  .GO(mid1_go), .port_62cc3b53_(bus_69808cf7_), .port_40cc1825_(bus_5ad36c45_), 
  .port_4c206d95_(bus_5122026c_), .port_4adb7c84_(bus_5122026c_), .port_7227ec97_(bus_52935bd9_), 
  .port_5277083b_(In1_DATA), .DONE(LL1_H_iunzipFilter2D_mid1_instance_DONE), 
  .RESULT(mid1), .RESULT_u98(mid1_u0), .RESULT_u99(mid1_u1), .RESULT_u100(mid1_u2), 
  .RESULT_u101(mid1_u3), .RESULT_u102(mid1_u4), .RESULT_u106(mid1_u5), .RESULT_u107(mid1_u6), 
  .RESULT_u108(mid1_u7), .RESULT_u109(mid1_u8), .RESULT_u103(mid1_u9), .RESULT_u104(mid1_u10), 
  .RESULT_u105(mid1_u11), .RESULT_u110(mid1_u12), .RESULT_u111(mid1_u13), .RESULT_u112(mid1_u14), 
  .RESULT_u113(mid1_u15));
LL1_H_iunzipFilter2D_midLeftNoConsume2 LL1_H_iunzipFilter2D_midLeftNoConsume2_instance(.CLK(CLK), 
  .RESET(bus_23506230_), .GO(midLeftNoConsume2_go), .port_5e0e4477_(16'h0), .port_11658ab7_(bus_5ad36c45_), 
  .port_77e7348e_(bus_78fb14d7_), .port_404d1402_(bus_27d78a2b_), .DONE(LL1_H_iunzipFilter2D_midLeftNoConsume2_instance_DONE), 
  .RESULT(midLeftNoConsume2), .RESULT_u114(midLeftNoConsume2_u0), .RESULT_u115(midLeftNoConsume2_u1), 
  .RESULT_u116(midLeftNoConsume2_u2), .RESULT_u117(midLeftNoConsume2_u3), .RESULT_u118(midLeftNoConsume2_u4), 
  .RESULT_u119(midLeftNoConsume2_u5), .RESULT_u120(midLeftNoConsume2_u6), .RESULT_u121(midLeftNoConsume2_u7), 
  .RESULT_u122(midLeftNoConsume2_u8));
assign bus_1564633b_=LL1_H_iunzipFilter2D_bottomRowNoConsume2_instance_DONE&{1{LL1_H_iunzipFilter2D_bottomRowNoConsume2_instance_DONE}};
LL1_H_iunzipFilter2D_stateVar_midPtr LL1_H_iunzipFilter2D_stateVar_midPtr_1(.bus_3400e46f_(CLK), 
  .bus_7a165d5a_(bus_23506230_), .bus_538c7874_(topLeft_u3), .bus_28a8a022_(topLeft_u4), 
  .bus_7badf2be_(topRow_u3), .bus_101c6579_(topRow_u4), .bus_5c59d90c_(topRight_u3), 
  .bus_1161e5a4_(16'h0), .bus_64256bdd_(midLeft1_u3), .bus_330204f5_(midLeft1_u4), 
  .bus_38b992ab_(midLeft2_u3), .bus_32076783_(midLeft2_u4), .bus_5a6e6bb4_(midLeftNoConsume1_u1), 
  .bus_4d247641_(midLeftNoConsume1_u2), .bus_7ed2fb60_(midLeftNoConsume2_u1), 
  .bus_65180804_(midLeftNoConsume2_u2), .bus_1be8c6a2_(mid1_u3), .bus_32f3848c_(mid1_u4), 
  .bus_5c9b2897_(mid2_u3), .bus_123ed54b_(mid2_u4), .bus_4f392724_(midNoConsume1_u1), 
  .bus_28004d89_(midNoConsume1_u2), .bus_7f3f31fb_(midNoConsume2_u1), .bus_1ba98a29_(midNoConsume2_u2), 
  .bus_2d59721d_(midRight1_u5), .bus_347ba71a_(16'h0), .bus_001a5c18_(midRight2_u5), 
  .bus_2eaf6154_(16'h0), .bus_32667a0e_(midRightNoConsume1_u1), .bus_0a10ed77_(16'h0), 
  .bus_1bfd9163_(midRightNoConsume2_u1), .bus_4d20b648_(16'h0), .bus_7151a5ac_(bottomLeftNoConsume1_u1), 
  .bus_4daa9a66_(bottomLeftNoConsume1_u2), .bus_35aa0d29_(bottomLeftNoConsume2_u1), 
  .bus_2ecb039d_(bottomLeftNoConsume2_u2), .bus_5730d21a_(bottomRowNoConsume1_u1), 
  .bus_48668b00_(bottomRowNoConsume1_u2), .bus_1910cc4e_(bottomRowNoConsume2_u1), 
  .bus_6613fb43_(bottomRowNoConsume2_u2), .bus_3ae651af_(bottomRightNoConsume1_u3), 
  .bus_53fb8955_(16'h0), .bus_2235ebf1_(bottomRightNoConsume2_u3), .bus_5a82cd0e_(16'h0), 
  .bus_5ad36c45_(bus_5ad36c45_));
assign bus_7a837774_=LL1_H_iunzipFilter2D_bottomLeftNoConsume1_instance_DONE&{1{LL1_H_iunzipFilter2D_bottomLeftNoConsume1_instance_DONE}};
assign bus_15ecd674_=LL1_H_iunzipFilter2D_midRightNoConsume1_instance_DONE&{1{LL1_H_iunzipFilter2D_midRightNoConsume1_instance_DONE}};
assign or_396b3042_u0=populateBuffer_u7|topLeft_u12|topRow_u14|topRight_u16|midLeft1_u12|midLeft2_u12|mid1_u12|mid2_u12|midRight1_u16|midRight2_u16;
LL1_H_iunzipFilter2D_simplememoryreferee_50b1249c_ LL1_H_iunzipFilter2D_simplememoryreferee_50b1249c__1(.bus_3d99ccb2_(CLK), 
  .bus_4561f8d0_(bus_23506230_), .bus_699bc1b7_(bus_02cec1f3_), .bus_5bec3b7f_(bus_25361c61_), 
  .bus_66b004a1_(populateBuffer_u3), .bus_3c867f89_(populateBuffer_u5), .bus_188ca39b_(populateBuffer_u4), 
  .bus_315688d8_(3'h1), .bus_7d411a66_(bus_7d411a66_), .bus_2da7af10_(bus_2da7af10_), 
  .bus_624df4b1_(bus_624df4b1_), .bus_3fffd7cb_(bus_3fffd7cb_), .bus_77051f23_(bus_77051f23_), 
  .bus_3681a366_(bus_3681a366_));
LL1_H_iunzipFilter2D_midLeft1 LL1_H_iunzipFilter2D_midLeft1_instance(.CLK(CLK), 
  .RESET(bus_23506230_), .GO(midLeft1_go), .port_7c96fb9c_(16'h0), .port_193dec0c_(bus_69808cf7_), 
  .port_3a87bf5f_(bus_5ad36c45_), .port_13cf03ae_(bus_7e378a50_), .port_76f10329_(bus_7e378a50_), 
  .port_32ad3201_(bus_167da5bd_), .port_718237b9_(In1_DATA), .DONE(LL1_H_iunzipFilter2D_midLeft1_instance_DONE), 
  .RESULT(midLeft1), .RESULT_u123(midLeft1_u0), .RESULT_u124(midLeft1_u1), .RESULT_u125(midLeft1_u2), 
  .RESULT_u126(midLeft1_u3), .RESULT_u127(midLeft1_u4), .RESULT_u131(midLeft1_u5), 
  .RESULT_u132(midLeft1_u6), .RESULT_u133(midLeft1_u7), .RESULT_u134(midLeft1_u8), 
  .RESULT_u128(midLeft1_u9), .RESULT_u129(midLeft1_u10), .RESULT_u130(midLeft1_u11), 
  .RESULT_u135(midLeft1_u12), .RESULT_u136(midLeft1_u13), .RESULT_u137(midLeft1_u14), 
  .RESULT_u138(midLeft1_u15));
assign bus_0379aee9_=LL1_H_iunzipFilter2D_midLeftNoConsume2_instance_DONE&{1{LL1_H_iunzipFilter2D_midLeftNoConsume2_instance_DONE}};
assign bus_73d09570_=LL1_H_iunzipFilter2D_midLeftNoConsume1_instance_DONE&{1{LL1_H_iunzipFilter2D_midLeftNoConsume1_instance_DONE}};
LL1_H_iunzipFilter2D_Kicker_6 LL1_H_iunzipFilter2D_Kicker_6_1(.CLK(CLK), .RESET(bus_23506230_), 
  .bus_4ae3b466_(bus_4ae3b466_));
assign or_0823cb19_u0=midLeft2_u14|midLeftNoConsume2_u7|mid2_u15|midNoConsume2_u8|midRight2_u18|midRightNoConsume2_u10|bottomLeftNoConsume2_u7|bottomRowNoConsume2_u8|bottomRightNoConsume2_u13;
assign bus_52c37c26_=LL1_H_iunzipFilter2D_topRight_instance_DONE&{1{LL1_H_iunzipFilter2D_topRight_instance_DONE}};
assign bus_46448f94_=LL1_H_iunzipFilter2D_donePopulateBuffer_instance_DONE&{1{LL1_H_iunzipFilter2D_donePopulateBuffer_instance_DONE}};
assign bus_12ce21da_=LL1_H_iunzipFilter2D_midRightNoConsume2_instance_DONE&{1{LL1_H_iunzipFilter2D_midRightNoConsume2_instance_DONE}};
assign bus_5d6bea1c_=LL1_H_iunzipFilter2D_mid1_instance_DONE&{1{LL1_H_iunzipFilter2D_mid1_instance_DONE}};
assign bus_4f3a32a9_=LL1_H_iunzipFilter2D_mid2_instance_DONE&{1{LL1_H_iunzipFilter2D_mid2_instance_DONE}};
LL1_H_iunzipFilter2D_donePopulateBuffer LL1_H_iunzipFilter2D_donePopulateBuffer_instance(.CLK(CLK), 
  .RESET(bus_23506230_), .GO(donePopulateBuffer_go), .DONE(LL1_H_iunzipFilter2D_donePopulateBuffer_instance_DONE), 
  .RESULT(donePopulateBuffer), .RESULT_u139(donePopulateBuffer_u0));
LL1_H_iunzipFilter2D_stateVar_fsmState_LL1_H_iunzipFilter2D LL1_H_iunzipFilter2D_stateVar_fsmState_LL1_H_iunzipFilter2D_1(.bus_3aa33e9e_(CLK), 
  .bus_0f971a50_(bus_23506230_), .bus_760e0512_(scheduler), .bus_628847e6_(scheduler_u18), 
  .bus_60d84d20_(bus_60d84d20_));
assign or_76a627f2_u0=midLeft2_u13|midLeftNoConsume2_u6|mid2_u13|midNoConsume2_u6|midRight2_u17|midRightNoConsume2_u8|bottomLeftNoConsume2_u6|bottomRowNoConsume2_u6|bottomRightNoConsume2_u12;
assign bus_4ca9c49f_=LL1_H_iunzipFilter2D_bottomLeftNoConsume2_instance_DONE&{1{LL1_H_iunzipFilter2D_bottomLeftNoConsume2_instance_DONE}};
LL1_H_iunzipFilter2D_bottomRightNoConsume1 LL1_H_iunzipFilter2D_bottomRightNoConsume1_instance(.CLK(CLK), 
  .RESET(bus_23506230_), .GO(bottomRightNoConsume1_go), .port_31e3635b_(bus_15ebb497_), 
  .port_43d1b2b6_(bus_6341aa95_), .port_4d9c680b_(bus_13a61289_), .DONE(LL1_H_iunzipFilter2D_bottomRightNoConsume1_instance_DONE), 
  .RESULT(bottomRightNoConsume1), .RESULT_u140(bottomRightNoConsume1_u0), .RESULT_u141(bottomRightNoConsume1_u1), 
  .RESULT_u142(bottomRightNoConsume1_u2), .RESULT_u143(bottomRightNoConsume1_u3), 
  .RESULT_u144(bottomRightNoConsume1_u4), .RESULT_u145(bottomRightNoConsume1_u5), 
  .RESULT_u146(bottomRightNoConsume1_u6), .RESULT_u147(bottomRightNoConsume1_u7), 
  .RESULT_u148(bottomRightNoConsume1_u8), .RESULT_u149(bottomRightNoConsume1_u9), 
  .RESULT_u150(bottomRightNoConsume1_u10), .RESULT_u151(bottomRightNoConsume1_u11), 
  .RESULT_u152(bottomRightNoConsume1_u12), .RESULT_u153(bottomRightNoConsume1_u13), 
  .RESULT_u154(bottomRightNoConsume1_u14));
LL1_H_iunzipFilter2D_stateVar_isEven LL1_H_iunzipFilter2D_stateVar_isEven_1(.bus_16c94a5f_(CLK), 
  .bus_06dd97a7_(bus_23506230_), .bus_23cf6553_(topRight_u7), .bus_1582983e_(topRight_u8), 
  .bus_193ba992_(midRight1_u7), .bus_250aabcd_(midRight1_u8), .bus_1503fca4_(midRight2_u7), 
  .bus_052f1bad_(midRight2_u8), .bus_5b66ba18_(midRightNoConsume1_u3), .bus_0fdbb770_(midRightNoConsume1_u4), 
  .bus_64dea1fa_(midRightNoConsume2_u3), .bus_652c6729_(midRightNoConsume2_u4), 
  .bus_4d350cfd_(bottomRightNoConsume1_u7), .bus_0dca5a75_(bottomRightNoConsume1_u8), 
  .bus_1946dfc4_(bottomRightNoConsume2_u7), .bus_06915c78_(bottomRightNoConsume2_u8), 
  .bus_15ebb497_(bus_15ebb497_));
LL1_H_iunzipFilter2D_bottomLeftNoConsume2 LL1_H_iunzipFilter2D_bottomLeftNoConsume2_instance(.CLK(CLK), 
  .RESET(bus_23506230_), .GO(bottomLeftNoConsume2_go), .port_773c7b8d_(16'h0), 
  .port_18be374b_(bus_5ad36c45_), .port_373fd3b4_(bus_0fd98caa_), .port_59b7d69f_(bus_623e353f_), 
  .DONE(LL1_H_iunzipFilter2D_bottomLeftNoConsume2_instance_DONE), .RESULT(bottomLeftNoConsume2), 
  .RESULT_u155(bottomLeftNoConsume2_u0), .RESULT_u156(bottomLeftNoConsume2_u1), 
  .RESULT_u157(bottomLeftNoConsume2_u2), .RESULT_u158(bottomLeftNoConsume2_u3), 
  .RESULT_u159(bottomLeftNoConsume2_u4), .RESULT_u160(bottomLeftNoConsume2_u5), 
  .RESULT_u161(bottomLeftNoConsume2_u6), .RESULT_u162(bottomLeftNoConsume2_u7), 
  .RESULT_u163(bottomLeftNoConsume2_u8));
LL1_H_iunzipFilter2D_topLeft LL1_H_iunzipFilter2D_topLeft_instance(.CLK(CLK), 
  .RESET(bus_23506230_), .GO(topLeft_go), .port_5221a8c5_(16'h0), .port_2026972c_(bus_69808cf7_), 
  .port_6d155da5_(bus_5ad36c45_), .port_792b0e97_(bus_295fc32e_), .port_20f4db23_(bus_7b6d2db0_), 
  .port_50f97c55_(bus_295fc32e_), .port_6e419463_(In1_DATA), .DONE(LL1_H_iunzipFilter2D_topLeft_instance_DONE), 
  .RESULT(topLeft), .RESULT_u164(topLeft_u0), .RESULT_u165(topLeft_u1), .RESULT_u166(topLeft_u2), 
  .RESULT_u167(topLeft_u3), .RESULT_u168(topLeft_u4), .RESULT_u169(topLeft_u5), 
  .RESULT_u170(topLeft_u6), .RESULT_u171(topLeft_u7), .RESULT_u172(topLeft_u8), 
  .RESULT_u173(topLeft_u9), .RESULT_u174(topLeft_u10), .RESULT_u175(topLeft_u11), 
  .RESULT_u176(topLeft_u12), .RESULT_u177(topLeft_u13), .RESULT_u178(topLeft_u14), 
  .RESULT_u179(topLeft_u15));
LL1_H_iunzipFilter2D_topRight LL1_H_iunzipFilter2D_topRight_instance(.CLK(CLK), 
  .RESET(bus_23506230_), .GO(topRight_go), .port_21a33c82_(bus_69808cf7_), .port_1f205dca_(bus_15ebb497_), 
  .port_468f8c2d_(bus_782a49ae_), .port_05847a01_(bus_75b6e6aa_), .port_0a351222_(bus_782a49ae_), 
  .port_19cb6266_(In1_DATA), .DONE(LL1_H_iunzipFilter2D_topRight_instance_DONE), 
  .RESULT(topRight), .RESULT_u180(topRight_u0), .RESULT_u181(topRight_u1), .RESULT_u182(topRight_u2), 
  .RESULT_u183(topRight_u3), .RESULT_u184(topRight_u4), .RESULT_u185(topRight_u5), 
  .RESULT_u186(topRight_u6), .RESULT_u187(topRight_u7), .RESULT_u188(topRight_u8), 
  .RESULT_u189(topRight_u9), .RESULT_u190(topRight_u10), .RESULT_u191(topRight_u11), 
  .RESULT_u192(topRight_u12), .RESULT_u193(topRight_u13), .RESULT_u194(topRight_u14), 
  .RESULT_u195(topRight_u15), .RESULT_u196(topRight_u16), .RESULT_u197(topRight_u17), 
  .RESULT_u198(topRight_u18), .RESULT_u199(topRight_u19));
LL1_H_iunzipFilter2D_structuralmemory_7648df26_ LL1_H_iunzipFilter2D_structuralmemory_7648df26__1(.CLK_u0(CLK), 
  .bus_7be93387_(bus_23506230_), .bus_500680a1_(bus_2da7af10_), .bus_14ede39e_(3'h1), 
  .bus_6f816ba1_(bus_3fffd7cb_), .bus_06d1faa7_(bus_624df4b1_), .bus_2ac66d9a_(bus_7d411a66_), 
  .bus_4cb922b4_(bus_1446f926_), .bus_7077ea2b_(3'h1), .bus_2b14349a_(bus_1df60b90_), 
  .bus_6e848c4c_(bus_7b461753_), .bus_6da7b786_(bus_1807f3cd_), .bus_25361c61_(bus_25361c61_), 
  .bus_02cec1f3_(bus_02cec1f3_), .bus_6dd7c8fd_(bus_6dd7c8fd_), .bus_7faecdeb_(bus_7faecdeb_));
LL1_H_iunzipFilter2D_midNoConsume1 LL1_H_iunzipFilter2D_midNoConsume1_instance(.CLK(CLK), 
  .RESET(bus_23506230_), .GO(midNoConsume1_go), .port_45028bf7_(bus_5ad36c45_), 
  .port_6e1d3735_(bus_57083dd4_), .port_55325b56_(bus_7cd6911c_), .DONE(LL1_H_iunzipFilter2D_midNoConsume1_instance_DONE), 
  .RESULT(midNoConsume1), .RESULT_u200(midNoConsume1_u0), .RESULT_u201(midNoConsume1_u1), 
  .RESULT_u202(midNoConsume1_u2), .RESULT_u203(midNoConsume1_u3), .RESULT_u204(midNoConsume1_u4), 
  .RESULT_u205(midNoConsume1_u5), .RESULT_u206(midNoConsume1_u6), .RESULT_u207(midNoConsume1_u7), 
  .RESULT_u208(midNoConsume1_u8));
LL1_H_iunzipFilter2D_midNoConsume2 LL1_H_iunzipFilter2D_midNoConsume2_instance(.CLK(CLK), 
  .RESET(bus_23506230_), .GO(midNoConsume2_go), .port_50b9449e_(bus_5ad36c45_), 
  .port_645796b3_(bus_0ad99597_), .port_7c5db129_(bus_2f7aa6e4_), .DONE(LL1_H_iunzipFilter2D_midNoConsume2_instance_DONE), 
  .RESULT(midNoConsume2), .RESULT_u209(midNoConsume2_u0), .RESULT_u210(midNoConsume2_u1), 
  .RESULT_u211(midNoConsume2_u2), .RESULT_u212(midNoConsume2_u3), .RESULT_u213(midNoConsume2_u4), 
  .RESULT_u214(midNoConsume2_u5), .RESULT_u215(midNoConsume2_u6), .RESULT_u216(midNoConsume2_u7), 
  .RESULT_u217(midNoConsume2_u8));
assign bus_1f82e86b_=LL1_H_iunzipFilter2D_midNoConsume2_instance_DONE&{1{LL1_H_iunzipFilter2D_midNoConsume2_instance_DONE}};
assign or_0315d09f_u0=midLeft2_u15|midLeftNoConsume2_u8|mid2_u14|midNoConsume2_u7|midRight2_u19|midRightNoConsume2_u9|bottomLeftNoConsume2_u8|bottomRowNoConsume2_u7|bottomRightNoConsume2_u14;
assign bus_6f5c9bce_=LL1_H_iunzipFilter2D_topLeft_instance_DONE&{1{LL1_H_iunzipFilter2D_topLeft_instance_DONE}};
assign bus_386c7386_=LL1_H_iunzipFilter2D_midNoConsume1_instance_DONE&{1{LL1_H_iunzipFilter2D_midNoConsume1_instance_DONE}};
LL1_H_iunzipFilter2D_simplememoryreferee_6b7a23db_ LL1_H_iunzipFilter2D_simplememoryreferee_6b7a23db__1(.bus_5baae8ff_(CLK), 
  .bus_7653fefb_(bus_23506230_), .bus_341c19c0_(bus_7faecdeb_), .bus_31af2b27_(bus_6dd7c8fd_), 
  .bus_3c374e45_(topLeft_u5), .bus_6913617c_(topLeft_u8), .bus_2cde6fec_(topLeft_u10), 
  .bus_3374a16b_(topLeft_u9), .bus_19f443bd_(3'h1), .bus_1553ab35_(topRow_u7), 
  .bus_663891ac_(topRow_u10), .bus_15e55fff_(topRow_u12), .bus_0d5861d7_(32'h0), 
  .bus_53cfd8c7_(3'h1), .bus_597c15fe_(topRight_u9), .bus_5900c238_(topRight_u12), 
  .bus_524805ba_(topRight_u14), .bus_3a1a33d5_(32'h0), .bus_3c586cf4_(3'h1), .bus_3c30ecac_(midLeft1_u9), 
  .bus_572c858a_(midLeft1_u5), .bus_75f74205_(midLeft1_u7), .bus_38f192ff_(32'h0), 
  .bus_675a6465_(3'h1), .bus_4185e507_(midLeft2_u9), .bus_38250251_(midLeft2_u5), 
  .bus_03b2b05f_(midLeft2_u7), .bus_7654652b_(32'h0), .bus_51b62008_(3'h1), .bus_5930e896_(midLeftNoConsume1_u3), 
  .bus_182c3189_(32'h0), .bus_472d9480_(3'h1), .bus_1ec5415f_(midLeftNoConsume2_u3), 
  .bus_1291fb88_(32'h0), .bus_0a2e3320_(3'h1), .bus_72eea4ff_(mid1_u9), .bus_77976b59_(mid1_u5), 
  .bus_3af85b4e_(mid1_u7), .bus_499884d1_(32'h0), .bus_1b25f6ba_(3'h1), .bus_74cb0e55_(mid2_u9), 
  .bus_756e636f_(mid2_u5), .bus_06803267_(mid2_u7), .bus_02376507_(32'h0), .bus_3be386e2_(3'h1), 
  .bus_013e7d74_(midNoConsume1_u3), .bus_37e5e149_(32'h0), .bus_0512548f_(3'h1), 
  .bus_398aca9c_(midNoConsume2_u3), .bus_007ee040_(32'h0), .bus_1d49e0c0_(3'h1), 
  .bus_1c6c6256_(midRight1_u13), .bus_08b6bf94_(midRight1_u9), .bus_06d6df27_(midRight1_u11), 
  .bus_74b6e615_(32'h0), .bus_63d1ee63_(3'h1), .bus_2a8034ec_(midRight2_u9), .bus_597f939d_(midRight2_u12), 
  .bus_309722e6_(midRight2_u14), .bus_783c1160_(32'h0), .bus_3295fff5_(3'h1), .bus_66b8fa73_(midRightNoConsume1_u5), 
  .bus_27bf1f93_(32'h0), .bus_56c466b1_(3'h1), .bus_3ab47106_(midRightNoConsume2_u5), 
  .bus_562d02e1_(32'h0), .bus_194c7c11_(3'h1), .bus_68a5f92c_(bottomLeftNoConsume1_u3), 
  .bus_3fe7f593_(32'h0), .bus_3c0153f0_(3'h1), .bus_22677e1d_(bottomLeftNoConsume2_u3), 
  .bus_0fc79387_(32'h0), .bus_55cc71ee_(3'h1), .bus_084108ff_(bottomRowNoConsume1_u3), 
  .bus_60937d22_(32'h0), .bus_39138d0a_(3'h1), .bus_38f0c907_(bottomRowNoConsume2_u3), 
  .bus_1be8460e_(32'h0), .bus_546e4ea1_(3'h1), .bus_68c80959_(bottomRightNoConsume1_u9), 
  .bus_723f4da1_(32'h0), .bus_118dcb12_(3'h1), .bus_34e6dfec_(bottomRightNoConsume2_u9), 
  .bus_47803ec7_(32'h0), .bus_5eb5ed16_(3'h1), .bus_1807f3cd_(bus_1807f3cd_), .bus_1446f926_(bus_1446f926_), 
  .bus_7b461753_(bus_7b461753_), .bus_1df60b90_(bus_1df60b90_), .bus_4ad1a98a_(bus_4ad1a98a_), 
  .bus_7b6d2db0_(bus_7b6d2db0_), .bus_295fc32e_(bus_295fc32e_), .bus_42424c02_(bus_42424c02_), 
  .bus_05553665_(bus_05553665_), .bus_75b6e6aa_(bus_75b6e6aa_), .bus_782a49ae_(bus_782a49ae_), 
  .bus_167da5bd_(bus_167da5bd_), .bus_7e378a50_(bus_7e378a50_), .bus_03a2926d_(bus_03a2926d_), 
  .bus_299c5c34_(bus_299c5c34_), .bus_12066278_(bus_12066278_), .bus_31710b5f_(bus_31710b5f_), 
  .bus_27d78a2b_(bus_27d78a2b_), .bus_78fb14d7_(bus_78fb14d7_), .bus_52935bd9_(bus_52935bd9_), 
  .bus_5122026c_(bus_5122026c_), .bus_35bb43c2_(bus_35bb43c2_), .bus_1f5c5926_(bus_1f5c5926_), 
  .bus_7cd6911c_(bus_7cd6911c_), .bus_57083dd4_(bus_57083dd4_), .bus_2f7aa6e4_(bus_2f7aa6e4_), 
  .bus_0ad99597_(bus_0ad99597_), .bus_5a5f2961_(bus_5a5f2961_), .bus_2781fc25_(bus_2781fc25_), 
  .bus_02c8854d_(bus_02c8854d_), .bus_3b77c854_(bus_3b77c854_), .bus_6308ab98_(bus_6308ab98_), 
  .bus_78addd53_(bus_78addd53_), .bus_2c656446_(bus_2c656446_), .bus_15fa8b31_(bus_15fa8b31_), 
  .bus_29c7540a_(bus_29c7540a_), .bus_24ac86a8_(bus_24ac86a8_), .bus_623e353f_(bus_623e353f_), 
  .bus_0fd98caa_(bus_0fd98caa_), .bus_4b3e6981_(bus_4b3e6981_), .bus_75734968_(bus_75734968_), 
  .bus_5727ff78_(bus_5727ff78_), .bus_018f435a_(bus_018f435a_), .bus_13a61289_(bus_13a61289_), 
  .bus_6341aa95_(bus_6341aa95_), .bus_5a1ddee7_(bus_5a1ddee7_), .bus_47b6d4cf_(bus_47b6d4cf_));
LL1_H_iunzipFilter2D_topRow LL1_H_iunzipFilter2D_topRow_instance(.CLK(CLK), .RESET(bus_23506230_), 
  .GO(topRow_go), .port_72b95caa_(bus_69808cf7_), .port_43ed3c0e_(bus_5ad36c45_), 
  .port_3b2ce771_(bus_4cb9b263_), .port_758e77d7_(bus_05553665_), .port_0b4ae4bc_(bus_42424c02_), 
  .port_59b37350_(bus_05553665_), .port_054c182e_(In1_DATA), .DONE(LL1_H_iunzipFilter2D_topRow_instance_DONE), 
  .RESULT(topRow), .RESULT_u218(topRow_u0), .RESULT_u219(topRow_u1), .RESULT_u220(topRow_u2), 
  .RESULT_u221(topRow_u3), .RESULT_u222(topRow_u4), .RESULT_u223(topRow_u5), .RESULT_u224(topRow_u6), 
  .RESULT_u225(topRow_u7), .RESULT_u226(topRow_u8), .RESULT_u227(topRow_u9), .RESULT_u228(topRow_u10), 
  .RESULT_u229(topRow_u11), .RESULT_u230(topRow_u12), .RESULT_u231(topRow_u13), 
  .RESULT_u232(topRow_u14), .RESULT_u233(topRow_u15), .RESULT_u234(topRow_u16), 
  .RESULT_u235(topRow_u17));
LL1_H_iunzipFilter2D_stateVar_idx LL1_H_iunzipFilter2D_stateVar_idx_1(.bus_0cf2d3f5_(CLK), 
  .bus_068d6c06_(bus_23506230_), .bus_674bf37e_(topLeft), .bus_10bc57e4_(16'h0), 
  .bus_4a2d20e1_(topRow_u1), .bus_22b29207_(16'h0), .bus_5c4dede9_(topRight_u1), 
  .bus_253147b9_(16'h0), .bus_4ebaa98e_(midLeft1), .bus_5ceaaebb_(16'h0), .bus_63833c02_(midLeft2), 
  .bus_50790775_(16'h0), .bus_2264995f_(midLeftNoConsume1), .bus_1cdbfe01_(16'h0), 
  .bus_2c539ca8_(midLeftNoConsume2), .bus_632c90cd_(16'h0), .bus_2397b779_(mid1_u1), 
  .bus_26b5b1f6_(16'h0), .bus_2570bc16_(mid2_u1), .bus_48005bbe_(16'h0), .bus_441deb71_(midNoConsume1), 
  .bus_46b2645c_(16'h0), .bus_62a23944_(midNoConsume2), .bus_1378e939_(16'h0), 
  .bus_513697cc_(midRight1), .bus_2cee4380_(16'h0), .bus_0475cc13_(midRight2), 
  .bus_78940204_(16'h0), .bus_766fd037_(bottomLeftNoConsume1), .bus_4d505dca_(16'h0), 
  .bus_1de90dae_(bottomLeftNoConsume2), .bus_20ace7e3_(16'h0), .bus_1c515fcc_(bottomRowNoConsume1), 
  .bus_5e13118c_(16'h0), .bus_041f2681_(bottomRowNoConsume2), .bus_6056c028_(16'h0), 
  .bus_3aa04241_(bottomRightNoConsume1_u1), .bus_3321cb07_(16'h0), .bus_7e50ec6c_(bottomRightNoConsume2_u1), 
  .bus_26d18263_(16'h0), .bus_2a7d4abb_(bus_2a7d4abb_));
LL1_H_iunzipFilter2D_midRight2 LL1_H_iunzipFilter2D_midRight2_instance(.CLK(CLK), 
  .RESET(bus_23506230_), .GO(midRight2_go), .port_5ef6bce8_(bus_69808cf7_), .port_5d219e2c_(bus_4cb9b263_), 
  .port_7888f833_(bus_15ebb497_), .port_0faf4797_(bus_3b77c854_), .port_46e25d42_(bus_02c8854d_), 
  .port_5cd1a04c_(bus_3b77c854_), .port_06fd2eaf_(In1_DATA), .DONE(LL1_H_iunzipFilter2D_midRight2_instance_DONE), 
  .RESULT(midRight2), .RESULT_u236(midRight2_u0), .RESULT_u237(midRight2_u1), .RESULT_u238(midRight2_u2), 
  .RESULT_u239(midRight2_u3), .RESULT_u240(midRight2_u4), .RESULT_u241(midRight2_u5), 
  .RESULT_u242(midRight2_u6), .RESULT_u243(midRight2_u7), .RESULT_u244(midRight2_u8), 
  .RESULT_u245(midRight2_u9), .RESULT_u246(midRight2_u10), .RESULT_u247(midRight2_u11), 
  .RESULT_u248(midRight2_u12), .RESULT_u249(midRight2_u13), .RESULT_u250(midRight2_u14), 
  .RESULT_u251(midRight2_u15), .RESULT_u252(midRight2_u16), .RESULT_u253(midRight2_u17), 
  .RESULT_u254(midRight2_u18), .RESULT_u255(midRight2_u19));
assign or_31aa5212_u0=topLeft_u15|topRow_u17|topRight_u19|midLeft1_u15|midLeftNoConsume1_u8|mid1_u15|midNoConsume1_u8|midRight1_u19|midRightNoConsume1_u10|bottomLeftNoConsume1_u8|bottomRowNoConsume1_u8|bottomRightNoConsume1_u14;
LL1_H_iunzipFilter2D_globalreset_physical_1f6e1ed4_ LL1_H_iunzipFilter2D_globalreset_physical_1f6e1ed4__1(.bus_68f6b794_(CLK), 
  .bus_1df2d7fb_(RESET), .bus_23506230_(bus_23506230_));
assign or_71cb5f0a_u0=topLeft_u13|topRow_u15|topRight_u17|midLeft1_u13|midLeftNoConsume1_u6|mid1_u13|midNoConsume1_u6|midRight1_u17|midRightNoConsume1_u8|bottomLeftNoConsume1_u6|bottomRowNoConsume1_u6|bottomRightNoConsume1_u12;
LL1_H_iunzipFilter2D_stateVar_processedRows LL1_H_iunzipFilter2D_stateVar_processedRows_1(.bus_50bd0603_(CLK), 
  .bus_06976a41_(bus_23506230_), .bus_334b47c1_(topRow_u5), .bus_360674e9_(topRow_u6), 
  .bus_2a00d576_(topRight_u5), .bus_52b2c6ce_(16'h1), .bus_5ab10369_(midRight1_u3), 
  .bus_7b0dad4e_(midRight1_u4), .bus_691edc7e_(midRight2_u3), .bus_2c378729_(midRight2_u4), 
  .bus_39e8dab6_(midRightNoConsume1), .bus_22ec21fb_(midRightNoConsume1_u0), 
  .bus_2bab2c65_(midRightNoConsume2), .bus_4dee9c66_(midRightNoConsume2_u0), 
  .bus_20abe20d_(bottomRightNoConsume1), .bus_6396d044_(16'h0), .bus_47b99ec4_(bottomRightNoConsume2), 
  .bus_5b45ada7_(16'h0), .bus_4cb9b263_(bus_4cb9b263_));
assign bus_67323e98_=LL1_H_iunzipFilter2D_midLeft1_instance_DONE&{1{LL1_H_iunzipFilter2D_midLeft1_instance_DONE}};
assign bus_6f12b7f2_=LL1_H_iunzipFilter2D_midLeft2_instance_DONE&{1{LL1_H_iunzipFilter2D_midLeft2_instance_DONE}};
LL1_H_iunzipFilter2D_bottomRightNoConsume2 LL1_H_iunzipFilter2D_bottomRightNoConsume2_instance(.CLK(CLK), 
  .RESET(bus_23506230_), .GO(bottomRightNoConsume2_go), .port_1379735b_(bus_15ebb497_), 
  .port_718e624c_(bus_47b6d4cf_), .port_680823aa_(bus_5a1ddee7_), .DONE(LL1_H_iunzipFilter2D_bottomRightNoConsume2_instance_DONE), 
  .RESULT(bottomRightNoConsume2), .RESULT_u256(bottomRightNoConsume2_u0), .RESULT_u257(bottomRightNoConsume2_u1), 
  .RESULT_u258(bottomRightNoConsume2_u2), .RESULT_u259(bottomRightNoConsume2_u3), 
  .RESULT_u260(bottomRightNoConsume2_u4), .RESULT_u261(bottomRightNoConsume2_u5), 
  .RESULT_u262(bottomRightNoConsume2_u6), .RESULT_u263(bottomRightNoConsume2_u7), 
  .RESULT_u264(bottomRightNoConsume2_u8), .RESULT_u265(bottomRightNoConsume2_u9), 
  .RESULT_u266(bottomRightNoConsume2_u10), .RESULT_u267(bottomRightNoConsume2_u11), 
  .RESULT_u268(bottomRightNoConsume2_u12), .RESULT_u269(bottomRightNoConsume2_u13), 
  .RESULT_u270(bottomRightNoConsume2_u14));
LL1_H_iunzipFilter2D_mid2 LL1_H_iunzipFilter2D_mid2_instance(.CLK(CLK), .RESET(bus_23506230_), 
  .GO(mid2_go), .port_63ca52d3_(bus_69808cf7_), .port_3ed342e9_(bus_5ad36c45_), 
  .port_22e17dd6_(bus_1f5c5926_), .port_61009e2d_(bus_1f5c5926_), .port_5174b1c2_(bus_35bb43c2_), 
  .port_28805c0d_(In1_DATA), .DONE(LL1_H_iunzipFilter2D_mid2_instance_DONE), 
  .RESULT(mid2), .RESULT_u271(mid2_u0), .RESULT_u272(mid2_u1), .RESULT_u273(mid2_u2), 
  .RESULT_u274(mid2_u3), .RESULT_u275(mid2_u4), .RESULT_u279(mid2_u5), .RESULT_u280(mid2_u6), 
  .RESULT_u281(mid2_u7), .RESULT_u282(mid2_u8), .RESULT_u276(mid2_u9), .RESULT_u277(mid2_u10), 
  .RESULT_u278(mid2_u11), .RESULT_u283(mid2_u12), .RESULT_u284(mid2_u13), .RESULT_u285(mid2_u14), 
  .RESULT_u286(mid2_u15));
LL1_H_iunzipFilter2D_bottomRowNoConsume2 LL1_H_iunzipFilter2D_bottomRowNoConsume2_instance(.CLK(CLK), 
  .RESET(bus_23506230_), .GO(bottomRowNoConsume2_go), .port_0c13a378_(bus_5ad36c45_), 
  .port_55afd2df_(bus_018f435a_), .port_137c836d_(bus_5727ff78_), .DONE(LL1_H_iunzipFilter2D_bottomRowNoConsume2_instance_DONE), 
  .RESULT(bottomRowNoConsume2), .RESULT_u287(bottomRowNoConsume2_u0), .RESULT_u288(bottomRowNoConsume2_u1), 
  .RESULT_u289(bottomRowNoConsume2_u2), .RESULT_u290(bottomRowNoConsume2_u3), 
  .RESULT_u291(bottomRowNoConsume2_u4), .RESULT_u292(bottomRowNoConsume2_u5), 
  .RESULT_u293(bottomRowNoConsume2_u6), .RESULT_u294(bottomRowNoConsume2_u7), 
  .RESULT_u295(bottomRowNoConsume2_u8));
assign bus_184376b1_=LL1_H_iunzipFilter2D_midRight1_instance_DONE&{1{LL1_H_iunzipFilter2D_midRight1_instance_DONE}};
assign or_4b5f8e83_u0=topLeft_u14|topRow_u16|topRight_u18|midLeft1_u14|midLeftNoConsume1_u7|mid1_u14|midNoConsume1_u7|midRight1_u18|midRightNoConsume1_u9|bottomLeftNoConsume1_u7|bottomRowNoConsume1_u7|bottomRightNoConsume1_u13;
assign bus_3fb35a7b_=LL1_H_iunzipFilter2D_bottomRightNoConsume2_instance_DONE&{1{LL1_H_iunzipFilter2D_bottomRightNoConsume2_instance_DONE}};
LL1_H_iunzipFilter2D_midLeft2 LL1_H_iunzipFilter2D_midLeft2_instance(.CLK(CLK), 
  .RESET(bus_23506230_), .GO(midLeft2_go), .port_55a161f7_(16'h0), .port_7ef80ea3_(bus_69808cf7_), 
  .port_0e0f96e7_(bus_5ad36c45_), .port_7b60df17_(bus_299c5c34_), .port_425dfc12_(bus_299c5c34_), 
  .port_1c2a9de3_(bus_03a2926d_), .port_17ab7fa3_(In1_DATA), .DONE(LL1_H_iunzipFilter2D_midLeft2_instance_DONE), 
  .RESULT(midLeft2), .RESULT_u296(midLeft2_u0), .RESULT_u297(midLeft2_u1), .RESULT_u298(midLeft2_u2), 
  .RESULT_u299(midLeft2_u3), .RESULT_u300(midLeft2_u4), .RESULT_u304(midLeft2_u5), 
  .RESULT_u305(midLeft2_u6), .RESULT_u306(midLeft2_u7), .RESULT_u307(midLeft2_u8), 
  .RESULT_u301(midLeft2_u9), .RESULT_u302(midLeft2_u10), .RESULT_u303(midLeft2_u11), 
  .RESULT_u308(midLeft2_u12), .RESULT_u309(midLeft2_u13), .RESULT_u310(midLeft2_u14), 
  .RESULT_u311(midLeft2_u15));
LL1_H_iunzipFilter2D_stateVar_consumed LL1_H_iunzipFilter2D_stateVar_consumed_1(.bus_29e3f084_(CLK), 
  .bus_3ddb8871_(bus_23506230_), .bus_41726d12_(populateBuffer_u1), .bus_16da44fd_(populateBuffer_u2), 
  .bus_742d05ab_(topLeft_u1), .bus_594dfb2b_(topLeft_u2), .bus_4c0950d8_(topRow), 
  .bus_4229c30d_(topRow_u0), .bus_3cf40804_(topRight), .bus_1b391612_(topRight_u0), 
  .bus_553e65f0_(midLeft1_u1), .bus_35213476_(midLeft1_u2), .bus_6df9cec0_(midLeft2_u1), 
  .bus_6e3ac2bf_(midLeft2_u2), .bus_777f8403_(mid1), .bus_3b684d2d_(mid1_u0), .bus_7ad94f9e_(mid2), 
  .bus_7a612d89_(mid2_u0), .bus_57752a3a_(midRight1_u1), .bus_6f16944e_(midRight1_u2), 
  .bus_77ad45a1_(midRight2_u1), .bus_7708085a_(midRight2_u2), .bus_5f8514a9_(bottomRightNoConsume1_u5), 
  .bus_7ee2b5b9_(32'h0), .bus_0da1a829_(bottomRightNoConsume2_u5), .bus_56da0d80_(32'h0), 
  .bus_69808cf7_(bus_69808cf7_));
LL1_H_iunzipFilter2D_stateVar_populatePtr LL1_H_iunzipFilter2D_stateVar_populatePtr_1(.bus_42988fd2_(CLK), 
  .bus_63643b3f_(bus_23506230_), .bus_65cf25d9_(populateBuffer), .bus_21d0a234_(populateBuffer_u0), 
  .bus_5fdc3a92_(donePopulateBuffer), .bus_668e6817_(16'h0), .bus_70eb3e5c_(bus_70eb3e5c_));
LL1_H_iunzipFilter2D_populateBuffer LL1_H_iunzipFilter2D_populateBuffer_instance(.CLK(CLK), 
  .RESET(bus_23506230_), .GO(populateBuffer_go), .port_623c9ece_(bus_70eb3e5c_), 
  .port_165a8581_(bus_69808cf7_), .port_7b608cd9_(bus_3681a366_), .port_4da138d8_(In1_DATA), 
  .DONE(LL1_H_iunzipFilter2D_populateBuffer_instance_DONE), .RESULT(populateBuffer), 
  .RESULT_u312(populateBuffer_u0), .RESULT_u313(populateBuffer_u1), .RESULT_u314(populateBuffer_u2), 
  .RESULT_u315(populateBuffer_u3), .RESULT_u316(populateBuffer_u4), .RESULT_u317(populateBuffer_u5), 
  .RESULT_u318(populateBuffer_u6), .RESULT_u319(populateBuffer_u7));
LL1_H_iunzipFilter2D_scheduler LL1_H_iunzipFilter2D_scheduler_instance(.CLK(CLK), 
  .RESET(bus_23506230_), .GO(bus_4ae3b466_), .port_42620ba7_(bus_60d84d20_), .port_41492b7c_(bus_70eb3e5c_), 
  .port_34f62b85_(bus_5ad36c45_), .port_6d2bfa2d_(bus_4cb9b263_), .port_2e0d86cd_(bus_69808cf7_), 
  .port_70e1f405_(bus_15ebb497_), .port_6d3af1f9_(In1_SEND), .port_459c8efa_(mid1_done), 
  .port_24157214_(bottomLeftNoConsume2_done), .port_6e290ca0_(midRight2_done), 
  .port_28187583_(bottomLeftNoConsume1_done), .port_5cc4abf1_(populateBuffer_done), 
  .port_010adde4_(bottomRightNoConsume2_done), .port_756b4eaa_(bottomRightNoConsume1_done), 
  .port_6004d831_(midRightNoConsume1_done), .port_0cc0d92d_(Out2_RDY), .port_4b42ea04_(bottomRowNoConsume1_done), 
  .port_6cf2bc2c_(topRow_done), .port_360d45ff_(midLeftNoConsume2_done), .port_213bddc2_(topLeft_done), 
  .port_0bf3d477_(midLeftNoConsume1_done), .port_24919790_(midRight1_done), .port_0cea4e99_(midLeft1_done), 
  .port_2374bcc1_(midLeft2_done), .port_1ff44368_(midNoConsume2_done), .port_1eaf7a9b_(mid2_done), 
  .port_40b0ff93_(topRight_done), .port_67286d84_(midNoConsume1_done), .port_4dcef735_(donePopulateBuffer_done), 
  .port_5e08959f_(Out1_RDY), .port_404885f8_(midRightNoConsume2_done), .port_6438f003_(bottomRowNoConsume2_done), 
  .DONE(LL1_H_iunzipFilter2D_scheduler_instance_DONE), .RESULT(scheduler), .RESULT_u320(scheduler_u18), 
  .RESULT_u321(scheduler_u19), .RESULT_u322(scheduler_u20), .RESULT_u323(scheduler_u21), 
  .RESULT_u324(scheduler_u22), .RESULT_u325(scheduler_u23), .RESULT_u326(scheduler_u24), 
  .RESULT_u327(scheduler_u25), .RESULT_u328(scheduler_u26), .RESULT_u329(scheduler_u27), 
  .RESULT_u330(scheduler_u28), .RESULT_u331(scheduler_u29), .RESULT_u332(scheduler_u30), 
  .RESULT_u333(scheduler_u31), .RESULT_u334(scheduler_u32), .RESULT_u335(scheduler_u33), 
  .RESULT_u336(scheduler_u34), .RESULT_u337(scheduler_u35), .RESULT_u338(scheduler_u36), 
  .RESULT_u339(scheduler_u37), .RESULT_u340(scheduler_u38), .RESULT_u341(scheduler_u39), 
  .RESULT_u342(scheduler_u40), .RESULT_u343(scheduler_u41));
LL1_H_iunzipFilter2D_midRightNoConsume1 LL1_H_iunzipFilter2D_midRightNoConsume1_instance(.CLK(CLK), 
  .RESET(bus_23506230_), .GO(midRightNoConsume1_go), .port_5a871a00_(bus_4cb9b263_), 
  .port_41319ec4_(bus_15ebb497_), .port_462e5940_(bus_78addd53_), .port_7baa5f0a_(bus_6308ab98_), 
  .DONE(LL1_H_iunzipFilter2D_midRightNoConsume1_instance_DONE), .RESULT(midRightNoConsume1), 
  .RESULT_u344(midRightNoConsume1_u0), .RESULT_u345(midRightNoConsume1_u1), .RESULT_u346(midRightNoConsume1_u2), 
  .RESULT_u347(midRightNoConsume1_u3), .RESULT_u348(midRightNoConsume1_u4), .RESULT_u349(midRightNoConsume1_u5), 
  .RESULT_u350(midRightNoConsume1_u6), .RESULT_u351(midRightNoConsume1_u7), .RESULT_u352(midRightNoConsume1_u8), 
  .RESULT_u353(midRightNoConsume1_u9), .RESULT_u354(midRightNoConsume1_u10));
assign bus_22299860_=LL1_H_iunzipFilter2D_midRight2_instance_DONE&{1{LL1_H_iunzipFilter2D_midRight2_instance_DONE}};
LL1_H_iunzipFilter2D_midRight1 LL1_H_iunzipFilter2D_midRight1_instance(.CLK(CLK), 
  .RESET(bus_23506230_), .GO(midRight1_go), .port_5330dddc_(bus_69808cf7_), .port_0e198730_(bus_4cb9b263_), 
  .port_55a91fbd_(bus_15ebb497_), .port_0ba14e5d_(bus_2781fc25_), .port_4d6b8630_(bus_2781fc25_), 
  .port_610b7aeb_(bus_5a5f2961_), .port_58e85b4e_(In1_DATA), .DONE(LL1_H_iunzipFilter2D_midRight1_instance_DONE), 
  .RESULT(midRight1), .RESULT_u355(midRight1_u0), .RESULT_u356(midRight1_u1), .RESULT_u357(midRight1_u2), 
  .RESULT_u358(midRight1_u3), .RESULT_u359(midRight1_u4), .RESULT_u360(midRight1_u5), 
  .RESULT_u361(midRight1_u6), .RESULT_u362(midRight1_u7), .RESULT_u363(midRight1_u8), 
  .RESULT_u367(midRight1_u9), .RESULT_u368(midRight1_u10), .RESULT_u369(midRight1_u11), 
  .RESULT_u370(midRight1_u12), .RESULT_u364(midRight1_u13), .RESULT_u365(midRight1_u14), 
  .RESULT_u366(midRight1_u15), .RESULT_u371(midRight1_u16), .RESULT_u372(midRight1_u17), 
  .RESULT_u373(midRight1_u18), .RESULT_u374(midRight1_u19));
endmodule



module LL1_H_iunzipFilter2D_midLeftNoConsume1(CLK, RESET, GO, port_24c1e388_, port_3d7d2b97_, port_4f846b64_, port_325dd0f8_, RESULT, RESULT_u60, RESULT_u61, RESULT_u62, RESULT_u63, RESULT_u64, RESULT_u65, RESULT_u66, RESULT_u67, RESULT_u68, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_24c1e388_;
input	[15:0]	port_3d7d2b97_;
input		port_4f846b64_;
input	[15:0]	port_325dd0f8_;
output		RESULT;
output	[15:0]	RESULT_u60;
output		RESULT_u61;
output	[15:0]	RESULT_u62;
output		RESULT_u63;
output	[31:0]	RESULT_u64;
output	[2:0]	RESULT_u65;
output	[15:0]	RESULT_u66;
output		RESULT_u67;
output	[15:0]	RESULT_u68;
output		DONE;
wire		or_u20_u0;
reg		done_cache_u0=1'h0;
wire		and_u104_u0;
reg		done_cache_u1_u0=1'h0;
wire		or_u21_u0;
wire		and_u109_u0;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_327e58bd_instance_RESULT;
wire	[15:0]	add;
wire		simplePinWrite;
wire	[15:0]	simplePinWrite_u28;
wire	[15:0]	simplePinWrite_u29;
reg		reg_2f819580_u0=1'h0;
reg		reg_00f1b5b4_u0=1'h0;
reg		reg_1bf7d58e_u0=1'h0;
reg		reg_1ac15051_u0=1'h0;
reg		reg_2f819580_result_delayed_u0=1'h0;
reg	[15:0]	syncEnable_u0=16'h0;
wire		or_u22_u0;
assign or_u20_u0=and_u104_u0|RESET;
always @(posedge CLK or posedge GO or posedge or_u20_u0)
begin
if (or_u20_u0)
done_cache_u0<=1'h0;
else if (GO)
done_cache_u0<=1'h1;
else done_cache_u0<=done_cache_u0;
end
assign and_u104_u0=done_cache_u0&port_4f846b64_;
always @(posedge CLK or posedge reg_1bf7d58e_u0 or posedge or_u21_u0)
begin
if (or_u21_u0)
done_cache_u1_u0<=1'h0;
else if (reg_1bf7d58e_u0)
done_cache_u1_u0<=1'h1;
else done_cache_u1_u0<=done_cache_u1_u0;
end
assign or_u21_u0=and_u109_u0|RESET;
assign and_u109_u0=done_cache_u1_u0&port_4f846b64_;
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_327e58bd_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_327e58bd_instance(.GO(reg_00f1b5b4_u0), 
  .port_1f5c7e5c_(syncEnable_u0), .port_01c233f0_(port_325dd0f8_), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_327e58bd_instance_RESULT));
assign add=port_3d7d2b97_+16'h1;
assign simplePinWrite=reg_00f1b5b4_u0&{1{reg_00f1b5b4_u0}};
assign simplePinWrite_u28=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_327e58bd_instance_RESULT&{16{reg_00f1b5b4_u0}};
assign simplePinWrite_u29=16'h1&{16{1'h1}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2f819580_u0<=1'h0;
else reg_2f819580_u0<=reg_00f1b5b4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00f1b5b4_u0<=1'h0;
else reg_00f1b5b4_u0<=reg_1bf7d58e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1bf7d58e_u0<=1'h0;
else reg_1bf7d58e_u0<=reg_1ac15051_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1ac15051_u0<=1'h0;
else reg_1ac15051_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2f819580_result_delayed_u0<=1'h0;
else reg_2f819580_result_delayed_u0<=reg_2f819580_u0;
end
always @(posedge CLK)
begin
if (reg_1ac15051_u0)
syncEnable_u0<=port_325dd0f8_;
end
assign or_u22_u0=GO|reg_1bf7d58e_u0;
assign RESULT=GO;
assign RESULT_u60=16'h0;
assign RESULT_u61=GO;
assign RESULT_u62=add;
assign RESULT_u63=or_u22_u0;
assign RESULT_u64=32'h0;
assign RESULT_u65=3'h1;
assign RESULT_u66=simplePinWrite_u29;
assign RESULT_u67=simplePinWrite;
assign RESULT_u68=simplePinWrite_u28;
assign DONE=reg_2f819580_result_delayed_u0;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_327e58bd_(GO, port_1f5c7e5c_, port_01c233f0_, RESULT);
input		GO;
input	[15:0]	port_1f5c7e5c_;
input	[15:0]	port_01c233f0_;
output	[15:0]	RESULT;
wire	[16:0]	add;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_1d4fe635_instance_RESULT;
assign add={port_1f5c7e5c_[15], port_1f5c7e5c_}+{port_01c233f0_[15], port_01c233f0_};
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_1d4fe635_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_1d4fe635_instance(.GO(GO), 
  .port_3d836049_({add[16], add[16:2]}), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_1d4fe635_instance_RESULT));
assign RESULT=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_1d4fe635_instance_RESULT;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_1d4fe635_(GO, port_3d836049_, RESULT);
input		GO;
input	[15:0]	port_3d836049_;
output	[15:0]	RESULT;
wire signed	[15:0]	greaterThan_a_signed;
wire signed	[15:0]	greaterThan_b_signed;
wire		greaterThan;
wire		and_u113_u0;
wire		and_u114_u0;
wire		not_u30_u0;
wire	[15:0]	mux_u8;
wire		and_u115_u0;
wire		and_u116_u0;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_3d836049_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign and_u113_u0=GO&not_u30_u0;
assign and_u114_u0=GO&greaterThan;
assign not_u30_u0=~greaterThan;
assign mux_u8=(and_u115_u0)?16'h0:port_3d836049_;
assign and_u115_u0=and_u114_u0&GO;
assign and_u116_u0=and_u113_u0&GO;
assign RESULT=mux_u8;
endmodule



module LL1_H_iunzipFilter2D_bottomRowNoConsume1(CLK, RESET, GO, port_72ef45b3_, port_6163a4df_, port_1df2cf41_, RESULT, RESULT_u69, RESULT_u70, RESULT_u71, RESULT_u72, RESULT_u73, RESULT_u74, RESULT_u75, RESULT_u76, RESULT_u77, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_72ef45b3_;
input		port_6163a4df_;
input	[15:0]	port_1df2cf41_;
output		RESULT;
output	[15:0]	RESULT_u69;
output		RESULT_u70;
output	[15:0]	RESULT_u71;
output		RESULT_u72;
output	[31:0]	RESULT_u73;
output	[2:0]	RESULT_u74;
output	[15:0]	RESULT_u75;
output		RESULT_u76;
output	[15:0]	RESULT_u77;
output		DONE;
wire		or_u23_u0;
reg		done_cache_u2=1'h0;
wire		and_u119_u0;
wire		or_u24_u0;
reg		done_cache_u3_u0=1'h0;
wire		and_u124_u0;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_495be67a_instance_RESULT;
wire	[15:0]	add;
wire	[15:0]	simplePinWrite;
wire	[15:0]	simplePinWrite_u30;
wire		simplePinWrite_u31;
reg		reg_7a084a03_u0=1'h0;
reg		reg_7141634e_u0=1'h0;
reg		reg_63060f4e_u0=1'h0;
reg		reg_7a084a03_result_delayed_u0=1'h0;
reg		reg_65deb06b_u0=1'h0;
wire		or_u25_u0;
reg	[15:0]	syncEnable_u1=16'h0;
assign or_u23_u0=and_u119_u0|RESET;
always @(posedge CLK or posedge GO or posedge or_u23_u0)
begin
if (or_u23_u0)
done_cache_u2<=1'h0;
else if (GO)
done_cache_u2<=1'h1;
else done_cache_u2<=done_cache_u2;
end
assign and_u119_u0=done_cache_u2&port_6163a4df_;
assign or_u24_u0=and_u124_u0|RESET;
always @(posedge CLK or posedge reg_7141634e_u0 or posedge or_u24_u0)
begin
if (or_u24_u0)
done_cache_u3_u0<=1'h0;
else if (reg_7141634e_u0)
done_cache_u3_u0<=1'h1;
else done_cache_u3_u0<=done_cache_u3_u0;
end
assign and_u124_u0=done_cache_u3_u0&port_6163a4df_;
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_495be67a_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_495be67a_instance(.GO(reg_7a084a03_u0), 
  .port_7447c3fa_(port_1df2cf41_), .port_61b39feb_(syncEnable_u1), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_495be67a_instance_RESULT));
assign add=port_72ef45b3_+16'h1;
assign simplePinWrite=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_495be67a_instance_RESULT&{16{reg_7a084a03_u0}};
assign simplePinWrite_u30=16'h1&{16{1'h1}};
assign simplePinWrite_u31=reg_7a084a03_u0&{1{reg_7a084a03_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a084a03_u0<=1'h0;
else reg_7a084a03_u0<=reg_7141634e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7141634e_u0<=1'h0;
else reg_7141634e_u0<=reg_65deb06b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_63060f4e_u0<=1'h0;
else reg_63060f4e_u0<=reg_7a084a03_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a084a03_result_delayed_u0<=1'h0;
else reg_7a084a03_result_delayed_u0<=reg_7a084a03_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_65deb06b_u0<=1'h0;
else reg_65deb06b_u0<=GO;
end
assign or_u25_u0=GO|reg_7141634e_u0;
always @(posedge CLK)
begin
if (reg_65deb06b_u0)
syncEnable_u1<=port_1df2cf41_;
end
assign RESULT=GO;
assign RESULT_u69=16'h0;
assign RESULT_u70=GO;
assign RESULT_u71=add;
assign RESULT_u72=or_u25_u0;
assign RESULT_u73=32'h0;
assign RESULT_u74=3'h1;
assign RESULT_u75=simplePinWrite_u30;
assign RESULT_u76=simplePinWrite_u31;
assign RESULT_u77=simplePinWrite;
assign DONE=reg_63060f4e_u0;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_495be67a_(GO, port_7447c3fa_, port_61b39feb_, RESULT);
input		GO;
input	[15:0]	port_7447c3fa_;
input	[15:0]	port_61b39feb_;
output	[15:0]	RESULT;
wire	[16:0]	add;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_44ab96d7_instance_RESULT;
assign add={port_61b39feb_[15], port_61b39feb_}+{port_7447c3fa_[15], port_7447c3fa_};
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_44ab96d7_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_44ab96d7_instance(.GO(GO), 
  .port_04e22c21_({add[16], add[16:2]}), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_44ab96d7_instance_RESULT));
assign RESULT=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_44ab96d7_instance_RESULT;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_44ab96d7_(GO, port_04e22c21_, RESULT);
input		GO;
input	[15:0]	port_04e22c21_;
output	[15:0]	RESULT;
wire signed	[15:0]	greaterThan_b_signed;
wire signed	[15:0]	greaterThan_a_signed;
wire		greaterThan;
wire		and_u128_u0;
wire		and_u129_u0;
wire		not_u31_u0;
wire	[15:0]	mux_u9;
wire		and_u130_u0;
wire		and_u131_u0;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_04e22c21_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign and_u128_u0=GO&not_u31_u0;
assign and_u129_u0=GO&greaterThan;
assign not_u31_u0=~greaterThan;
assign mux_u9=(and_u131_u0)?port_04e22c21_:16'h0;
assign and_u130_u0=and_u129_u0&GO;
assign and_u131_u0=and_u128_u0&GO;
assign RESULT=mux_u9;
endmodule



module LL1_H_iunzipFilter2D_midRightNoConsume2(CLK, RESET, GO, port_461847e8_, port_24a7300a_, port_03e1c37e_, port_0d8191ee_, RESULT, RESULT_u78, RESULT_u79, RESULT_u80, RESULT_u81, RESULT_u82, RESULT_u83, RESULT_u84, RESULT_u85, RESULT_u86, RESULT_u87, RESULT_u88, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_461847e8_;
input		port_24a7300a_;
input		port_03e1c37e_;
input	[15:0]	port_0d8191ee_;
output		RESULT;
output	[15:0]	RESULT_u78;
output		RESULT_u79;
output	[15:0]	RESULT_u80;
output		RESULT_u81;
output		RESULT_u82;
output		RESULT_u83;
output	[31:0]	RESULT_u84;
output	[2:0]	RESULT_u85;
output	[15:0]	RESULT_u86;
output	[15:0]	RESULT_u87;
output		RESULT_u88;
output		DONE;
reg		done_cache_u4=1'h0;
wire		or_u26_u0;
wire		and_u134_u0;
reg		done_cache_u5_u0=1'h0;
wire		or_u27_u0;
wire		and_u139_u0;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_06a80709_instance_RESULT;
wire	[15:0]	add;
wire		not_u33;
wire	[15:0]	simplePinWrite;
wire	[15:0]	simplePinWrite_u32;
wire		simplePinWrite_u33;
reg		reg_27ad8383_u0=1'h0;
reg		reg_6ac062a6_u0=1'h0;
reg		reg_33e42890_u0=1'h0;
reg		reg_629b351b_u0=1'h0;
reg		reg_27ad8383_result_delayed_u0=1'h0;
reg	[15:0]	syncEnable_u2=16'h0;
wire		or_u28_u0;
always @(posedge CLK or posedge GO or posedge or_u26_u0)
begin
if (or_u26_u0)
done_cache_u4<=1'h0;
else if (GO)
done_cache_u4<=1'h1;
else done_cache_u4<=done_cache_u4;
end
assign or_u26_u0=and_u134_u0|RESET;
assign and_u134_u0=done_cache_u4&port_03e1c37e_;
always @(posedge CLK or posedge reg_27ad8383_u0 or posedge or_u27_u0)
begin
if (or_u27_u0)
done_cache_u5_u0<=1'h0;
else if (reg_27ad8383_u0)
done_cache_u5_u0<=1'h1;
else done_cache_u5_u0<=done_cache_u5_u0;
end
assign or_u27_u0=and_u139_u0|RESET;
assign and_u139_u0=done_cache_u5_u0&port_03e1c37e_;
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_06a80709_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_06a80709_instance(.GO(reg_27ad8383_result_delayed_u0), 
  .port_4d0b894d_(syncEnable_u2), .port_665b6c28_(port_0d8191ee_), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_06a80709_instance_RESULT));
assign add=port_461847e8_+16'h1;
assign not_u33=!port_24a7300a_;
assign simplePinWrite=16'h1&{16{1'h1}};
assign simplePinWrite_u32=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_06a80709_instance_RESULT&{16{reg_27ad8383_result_delayed_u0}};
assign simplePinWrite_u33=reg_27ad8383_result_delayed_u0&{1{reg_27ad8383_result_delayed_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_27ad8383_u0<=1'h0;
else reg_27ad8383_u0<=reg_6ac062a6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6ac062a6_u0<=1'h0;
else reg_6ac062a6_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_33e42890_u0<=1'h0;
else reg_33e42890_u0<=reg_629b351b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_629b351b_u0<=1'h0;
else reg_629b351b_u0<=reg_27ad8383_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_27ad8383_result_delayed_u0<=1'h0;
else reg_27ad8383_result_delayed_u0<=reg_27ad8383_u0;
end
always @(posedge CLK)
begin
if (reg_6ac062a6_u0)
syncEnable_u2<=port_0d8191ee_;
end
assign or_u28_u0=GO|reg_27ad8383_u0;
assign RESULT=GO;
assign RESULT_u78=add;
assign RESULT_u79=GO;
assign RESULT_u80=16'h0;
assign RESULT_u81=GO;
assign RESULT_u82=not_u33;
assign RESULT_u83=or_u28_u0;
assign RESULT_u84=32'h0;
assign RESULT_u85=3'h1;
assign RESULT_u86=simplePinWrite;
assign RESULT_u87=simplePinWrite_u32;
assign RESULT_u88=simplePinWrite_u33;
assign DONE=reg_33e42890_u0;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_06a80709_(GO, port_4d0b894d_, port_665b6c28_, RESULT);
input		GO;
input	[15:0]	port_4d0b894d_;
input	[15:0]	port_665b6c28_;
output	[15:0]	RESULT;
wire	[15:0]	subtract;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_31df6d88_instance_RESULT;
assign subtract=port_4d0b894d_-port_665b6c28_;
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_31df6d88_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_31df6d88_instance(.GO(GO), 
  .port_0aab2900_({subtract[15], subtract[15:1]}), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_31df6d88_instance_RESULT));
assign RESULT=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_31df6d88_instance_RESULT;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_31df6d88_(GO, port_0aab2900_, RESULT);
input		GO;
input	[15:0]	port_0aab2900_;
output	[15:0]	RESULT;
wire signed	[15:0]	greaterThan_b_signed;
wire		greaterThan;
wire signed	[15:0]	greaterThan_a_signed;
wire		not_u32_u0;
wire		and_u143_u0;
wire		and_u144_u0;
wire		and_u145_u0;
wire		and_u146_u0;
wire	[15:0]	mux_u10;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_0aab2900_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign not_u32_u0=~greaterThan;
assign and_u143_u0=GO&not_u32_u0;
assign and_u144_u0=GO&greaterThan;
assign and_u145_u0=and_u144_u0&GO;
assign and_u146_u0=and_u143_u0&GO;
assign mux_u10=(and_u145_u0)?16'h0:port_0aab2900_;
assign RESULT=mux_u10;
endmodule



module LL1_H_iunzipFilter2D_bottomLeftNoConsume1(CLK, RESET, GO, port_47f3deda_, port_01459c00_, port_4b02a40f_, port_5e56587d_, RESULT, RESULT_u89, RESULT_u90, RESULT_u91, RESULT_u92, RESULT_u93, RESULT_u94, RESULT_u95, RESULT_u96, RESULT_u97, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_47f3deda_;
input	[15:0]	port_01459c00_;
input		port_4b02a40f_;
input	[15:0]	port_5e56587d_;
output		RESULT;
output	[15:0]	RESULT_u89;
output		RESULT_u90;
output	[15:0]	RESULT_u91;
output		RESULT_u92;
output	[31:0]	RESULT_u93;
output	[2:0]	RESULT_u94;
output	[15:0]	RESULT_u95;
output		RESULT_u96;
output	[15:0]	RESULT_u97;
output		DONE;
wire		and_u147_u0;
wire		or_u29_u0;
reg		done_cache_u6=1'h0;
reg		done_cache_u7_u0=1'h0;
wire		and_u152_u0;
wire		or_u30_u0;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_54fec8e2_instance_RESULT;
wire	[15:0]	add;
wire	[15:0]	simplePinWrite;
wire	[15:0]	simplePinWrite_u34;
wire		simplePinWrite_u35;
reg		reg_3efc0af3_u0=1'h0;
reg		reg_0b8d3393_u0=1'h0;
reg		reg_443dc122_u0=1'h0;
reg	[15:0]	syncEnable_u3=16'h0;
reg		reg_3efc0af3_result_delayed_u0=1'h0;
wire		or_u31_u0;
reg		reg_443dc122_result_delayed_u0=1'h0;
assign and_u147_u0=done_cache_u6&port_4b02a40f_;
assign or_u29_u0=and_u147_u0|RESET;
always @(posedge CLK or posedge GO or posedge or_u29_u0)
begin
if (or_u29_u0)
done_cache_u6<=1'h0;
else if (GO)
done_cache_u6<=1'h1;
else done_cache_u6<=done_cache_u6;
end
always @(posedge CLK or posedge reg_3efc0af3_result_delayed_u0 or posedge or_u30_u0)
begin
if (or_u30_u0)
done_cache_u7_u0<=1'h0;
else if (reg_3efc0af3_result_delayed_u0)
done_cache_u7_u0<=1'h1;
else done_cache_u7_u0<=done_cache_u7_u0;
end
assign and_u152_u0=done_cache_u7_u0&port_4b02a40f_;
assign or_u30_u0=and_u152_u0|RESET;
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_54fec8e2_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_54fec8e2_instance(.GO(reg_443dc122_u0), 
  .port_2589646e_(syncEnable_u3), .port_4084d7a9_(port_5e56587d_), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_54fec8e2_instance_RESULT));
assign add=port_01459c00_+16'h1;
assign simplePinWrite=16'h1&{16{1'h1}};
assign simplePinWrite_u34=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_54fec8e2_instance_RESULT&{16{reg_443dc122_u0}};
assign simplePinWrite_u35=reg_443dc122_u0&{1{reg_443dc122_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3efc0af3_u0<=1'h0;
else reg_3efc0af3_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0b8d3393_u0<=1'h0;
else reg_0b8d3393_u0<=reg_443dc122_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_443dc122_u0<=1'h0;
else reg_443dc122_u0<=reg_3efc0af3_result_delayed_u0;
end
always @(posedge CLK)
begin
if (reg_3efc0af3_u0)
syncEnable_u3<=port_5e56587d_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3efc0af3_result_delayed_u0<=1'h0;
else reg_3efc0af3_result_delayed_u0<=reg_3efc0af3_u0;
end
assign or_u31_u0=GO|reg_3efc0af3_result_delayed_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_443dc122_result_delayed_u0<=1'h0;
else reg_443dc122_result_delayed_u0<=reg_443dc122_u0;
end
assign RESULT=GO;
assign RESULT_u89=16'h0;
assign RESULT_u90=GO;
assign RESULT_u91=add;
assign RESULT_u92=or_u31_u0;
assign RESULT_u93=32'h0;
assign RESULT_u94=3'h1;
assign RESULT_u95=simplePinWrite;
assign RESULT_u96=simplePinWrite_u35;
assign RESULT_u97=simplePinWrite_u34;
assign DONE=reg_0b8d3393_u0;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_54fec8e2_(GO, port_2589646e_, port_4084d7a9_, RESULT);
input		GO;
input	[15:0]	port_2589646e_;
input	[15:0]	port_4084d7a9_;
output	[15:0]	RESULT;
wire	[16:0]	add;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_60c3fa96_instance_RESULT;
assign add={port_2589646e_[15], port_2589646e_}+{port_4084d7a9_[15], port_4084d7a9_};
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_60c3fa96_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_60c3fa96_instance(.GO(GO), 
  .port_14955648_({add[16], add[16:2]}), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_60c3fa96_instance_RESULT));
assign RESULT=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_60c3fa96_instance_RESULT;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_60c3fa96_(GO, port_14955648_, RESULT);
input		GO;
input	[15:0]	port_14955648_;
output	[15:0]	RESULT;
wire signed	[15:0]	greaterThan_b_signed;
wire		greaterThan;
wire signed	[15:0]	greaterThan_a_signed;
wire		and_u156_u0;
wire		and_u157_u0;
wire		not_u34_u0;
wire		and_u158_u0;
wire	[15:0]	mux_u11;
wire		and_u159_u0;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_14955648_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign and_u156_u0=GO&not_u34_u0;
assign and_u157_u0=GO&greaterThan;
assign not_u34_u0=~greaterThan;
assign and_u158_u0=and_u157_u0&GO;
assign mux_u11=(and_u158_u0)?16'h0:port_14955648_;
assign and_u159_u0=and_u156_u0&GO;
assign RESULT=mux_u11;
endmodule



module LL1_H_iunzipFilter2D_mid1(CLK, RESET, GO, port_62cc3b53_, port_40cc1825_, port_4adb7c84_, port_7227ec97_, port_4c206d95_, port_5277083b_, RESULT, RESULT_u98, RESULT_u99, RESULT_u100, RESULT_u101, RESULT_u102, RESULT_u103, RESULT_u104, RESULT_u105, RESULT_u106, RESULT_u107, RESULT_u108, RESULT_u109, RESULT_u110, RESULT_u111, RESULT_u112, RESULT_u113, DONE);
input		CLK;
input		RESET;
input		GO;
input	[31:0]	port_62cc3b53_;
input	[15:0]	port_40cc1825_;
input		port_4adb7c84_;
input	[15:0]	port_7227ec97_;
input		port_4c206d95_;
input	[15:0]	port_5277083b_;
output		RESULT;
output	[31:0]	RESULT_u98;
output		RESULT_u99;
output	[15:0]	RESULT_u100;
output		RESULT_u101;
output	[15:0]	RESULT_u102;
output		RESULT_u103;
output	[31:0]	RESULT_u104;
output	[2:0]	RESULT_u105;
output		RESULT_u106;
output	[31:0]	RESULT_u107;
output	[15:0]	RESULT_u108;
output	[2:0]	RESULT_u109;
output		RESULT_u110;
output	[15:0]	RESULT_u111;
output		RESULT_u112;
output	[15:0]	RESULT_u113;
output		DONE;
wire		simplePinWrite;
reg		done_cache_u8=1'h0;
wire		or_u32_u0;
wire		and_u162_u0;
reg		done_cache_u9_u0=1'h0;
wire		and_u167_u0;
wire		or_u33_u0;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_393aa8a3_instance_RESULT;
wire		and_u176_u0;
wire		or_u34_u0;
reg		reg_52cba022_u0=1'h0;
wire	[31:0]	add;
wire	[15:0]	add_u0;
wire		simplePinWrite_u36;
wire	[15:0]	simplePinWrite_u37;
wire	[15:0]	simplePinWrite_u38;
reg		reg_38acca9e_u0=1'h0;
reg		reg_56a8b09e_u0=1'h0;
reg	[15:0]	syncEnable_u4=16'h0;
reg	[15:0]	syncEnable_u5_u0=16'h0;
reg		reg_56a8b09e_result_delayed_u0=1'h0;
reg		reg_4846bd59_u0=1'h0;
reg		reg_56a8b09e_result_delayed_result_delayed_u0=1'h0;
wire		or_u35_u0;
reg		reg_38acca9e_result_delayed_u0=1'h0;
assign simplePinWrite=GO&{1{GO}};
always @(posedge CLK or posedge GO or posedge or_u32_u0)
begin
if (or_u32_u0)
done_cache_u8<=1'h0;
else if (GO)
done_cache_u8<=1'h1;
else done_cache_u8<=done_cache_u8;
end
assign or_u32_u0=and_u162_u0|RESET;
assign and_u162_u0=done_cache_u8&port_4c206d95_;
always @(posedge CLK or posedge reg_38acca9e_u0 or posedge or_u33_u0)
begin
if (or_u33_u0)
done_cache_u9_u0<=1'h0;
else if (reg_38acca9e_u0)
done_cache_u9_u0<=1'h1;
else done_cache_u9_u0<=done_cache_u9_u0;
end
assign and_u167_u0=done_cache_u9_u0&port_4c206d95_;
assign or_u33_u0=and_u167_u0|RESET;
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_393aa8a3_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_393aa8a3_instance(.GO(reg_38acca9e_result_delayed_u0), 
  .port_129098d2_(port_7227ec97_), .port_1b1a0f51_(syncEnable_u4), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_393aa8a3_instance_RESULT));
assign and_u176_u0=reg_52cba022_u0&port_4c206d95_;
assign or_u34_u0=and_u176_u0|RESET;
always @(posedge CLK or posedge reg_56a8b09e_result_delayed_u0 or posedge or_u34_u0)
begin
if (or_u34_u0)
reg_52cba022_u0<=1'h0;
else if (reg_56a8b09e_result_delayed_u0)
reg_52cba022_u0<=1'h1;
else reg_52cba022_u0<=reg_52cba022_u0;
end
assign add=port_62cc3b53_+32'h1;
assign add_u0=port_40cc1825_+16'h1;
assign simplePinWrite_u36=reg_38acca9e_result_delayed_u0&{1{reg_38acca9e_result_delayed_u0}};
assign simplePinWrite_u37=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_393aa8a3_instance_RESULT&{16{reg_38acca9e_result_delayed_u0}};
assign simplePinWrite_u38=16'h1&{16{1'h1}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_38acca9e_u0<=1'h0;
else reg_38acca9e_u0<=reg_4846bd59_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_56a8b09e_u0<=1'h0;
else reg_56a8b09e_u0<=reg_38acca9e_result_delayed_u0;
end
always @(posedge CLK)
begin
if (reg_4846bd59_u0)
syncEnable_u4<=port_7227ec97_;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u5_u0<=port_5277083b_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_56a8b09e_result_delayed_u0<=1'h0;
else reg_56a8b09e_result_delayed_u0<=reg_56a8b09e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4846bd59_u0<=1'h0;
else reg_4846bd59_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_56a8b09e_result_delayed_result_delayed_u0<=1'h0;
else reg_56a8b09e_result_delayed_result_delayed_u0<=reg_56a8b09e_result_delayed_u0;
end
assign or_u35_u0=GO|reg_38acca9e_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_38acca9e_result_delayed_u0<=1'h0;
else reg_38acca9e_result_delayed_u0<=reg_38acca9e_u0;
end
assign RESULT=GO;
assign RESULT_u98=add;
assign RESULT_u99=GO;
assign RESULT_u100=16'h0;
assign RESULT_u101=GO;
assign RESULT_u102=add_u0;
assign RESULT_u103=or_u35_u0;
assign RESULT_u104=32'h0;
assign RESULT_u105=3'h1;
assign RESULT_u106=reg_56a8b09e_result_delayed_u0;
assign RESULT_u107=32'h0;
assign RESULT_u108=syncEnable_u5_u0;
assign RESULT_u109=3'h1;
assign RESULT_u110=simplePinWrite;
assign RESULT_u111=simplePinWrite_u38;
assign RESULT_u112=simplePinWrite_u36;
assign RESULT_u113=simplePinWrite_u37;
assign DONE=reg_56a8b09e_result_delayed_result_delayed_u0;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_393aa8a3_(GO, port_129098d2_, port_1b1a0f51_, RESULT);
input		GO;
input	[15:0]	port_129098d2_;
input	[15:0]	port_1b1a0f51_;
output	[15:0]	RESULT;
wire	[16:0]	add;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_1761f8df_instance_RESULT;
assign add={port_1b1a0f51_[15], port_1b1a0f51_}+{port_129098d2_[15], port_129098d2_};
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_1761f8df_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_1761f8df_instance(.GO(GO), 
  .port_411d8326_({add[16], add[16:2]}), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_1761f8df_instance_RESULT));
assign RESULT=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_1761f8df_instance_RESULT;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_1761f8df_(GO, port_411d8326_, RESULT);
input		GO;
input	[15:0]	port_411d8326_;
output	[15:0]	RESULT;
wire signed	[15:0]	greaterThan_b_signed;
wire signed	[15:0]	greaterThan_a_signed;
wire		greaterThan;
wire		and_u171_u0;
wire		not_u35_u0;
wire		and_u172_u0;
wire		and_u173_u0;
wire		and_u174_u0;
wire	[15:0]	mux_u12;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_411d8326_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign and_u171_u0=GO&not_u35_u0;
assign not_u35_u0=~greaterThan;
assign and_u172_u0=GO&greaterThan;
assign and_u173_u0=and_u172_u0&GO;
assign and_u174_u0=and_u171_u0&GO;
assign mux_u12=(and_u173_u0)?16'h0:port_411d8326_;
assign RESULT=mux_u12;
endmodule



module LL1_H_iunzipFilter2D_midLeftNoConsume2(CLK, RESET, GO, port_5e0e4477_, port_11658ab7_, port_77e7348e_, port_404d1402_, RESULT, RESULT_u114, RESULT_u115, RESULT_u116, RESULT_u117, RESULT_u118, RESULT_u119, RESULT_u120, RESULT_u121, RESULT_u122, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_5e0e4477_;
input	[15:0]	port_11658ab7_;
input		port_77e7348e_;
input	[15:0]	port_404d1402_;
output		RESULT;
output	[15:0]	RESULT_u114;
output		RESULT_u115;
output	[15:0]	RESULT_u116;
output		RESULT_u117;
output	[31:0]	RESULT_u118;
output	[2:0]	RESULT_u119;
output	[15:0]	RESULT_u120;
output		RESULT_u121;
output	[15:0]	RESULT_u122;
output		DONE;
reg		done_cache_u10=1'h0;
wire		or_u36_u0;
wire		and_u178_u0;
reg		done_cache_u11_u0=1'h0;
wire		and_u183_u0;
wire		or_u37_u0;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_09e6e252_instance_RESULT;
wire	[15:0]	add;
wire	[15:0]	simplePinWrite;
wire		simplePinWrite_u39;
wire	[15:0]	simplePinWrite_u40;
reg		reg_49f0ded8_u0=1'h0;
wire		or_u38_u0;
reg	[15:0]	syncEnable_u6=16'h0;
reg		reg_44bded3c_u0=1'h0;
reg		reg_075acbde_u0=1'h0;
reg		reg_570f0cce_u0=1'h0;
reg		reg_44bded3c_result_delayed_u0=1'h0;
always @(posedge CLK or posedge GO or posedge or_u36_u0)
begin
if (or_u36_u0)
done_cache_u10<=1'h0;
else if (GO)
done_cache_u10<=1'h1;
else done_cache_u10<=done_cache_u10;
end
assign or_u36_u0=and_u178_u0|RESET;
assign and_u178_u0=done_cache_u10&port_77e7348e_;
always @(posedge CLK or posedge reg_44bded3c_u0 or posedge or_u37_u0)
begin
if (or_u37_u0)
done_cache_u11_u0<=1'h0;
else if (reg_44bded3c_u0)
done_cache_u11_u0<=1'h1;
else done_cache_u11_u0<=done_cache_u11_u0;
end
assign and_u183_u0=done_cache_u11_u0&port_77e7348e_;
assign or_u37_u0=and_u183_u0|RESET;
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_09e6e252_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_09e6e252_instance(.GO(reg_44bded3c_result_delayed_u0), 
  .port_2530552c_(syncEnable_u6), .port_7f37585b_(port_404d1402_), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_09e6e252_instance_RESULT));
assign add=port_11658ab7_+16'h1;
assign simplePinWrite=16'h1&{16{1'h1}};
assign simplePinWrite_u39=reg_44bded3c_result_delayed_u0&{1{reg_44bded3c_result_delayed_u0}};
assign simplePinWrite_u40=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_09e6e252_instance_RESULT&{16{reg_44bded3c_result_delayed_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_49f0ded8_u0<=1'h0;
else reg_49f0ded8_u0<=reg_570f0cce_u0;
end
assign or_u38_u0=GO|reg_44bded3c_u0;
always @(posedge CLK)
begin
if (reg_075acbde_u0)
syncEnable_u6<=port_404d1402_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_44bded3c_u0<=1'h0;
else reg_44bded3c_u0<=reg_075acbde_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_075acbde_u0<=1'h0;
else reg_075acbde_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_570f0cce_u0<=1'h0;
else reg_570f0cce_u0<=reg_44bded3c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_44bded3c_result_delayed_u0<=1'h0;
else reg_44bded3c_result_delayed_u0<=reg_44bded3c_u0;
end
assign RESULT=GO;
assign RESULT_u114=16'h0;
assign RESULT_u115=GO;
assign RESULT_u116=add;
assign RESULT_u117=or_u38_u0;
assign RESULT_u118=32'h0;
assign RESULT_u119=3'h1;
assign RESULT_u120=simplePinWrite;
assign RESULT_u121=simplePinWrite_u39;
assign RESULT_u122=simplePinWrite_u40;
assign DONE=reg_49f0ded8_u0;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_09e6e252_(GO, port_2530552c_, port_7f37585b_, RESULT);
input		GO;
input	[15:0]	port_2530552c_;
input	[15:0]	port_7f37585b_;
output	[15:0]	RESULT;
wire	[15:0]	subtract;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_40446f2e_instance_RESULT;
assign subtract=port_2530552c_-port_7f37585b_;
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_40446f2e_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_40446f2e_instance(.GO(GO), 
  .port_3bf115d5_({subtract[15], subtract[15:1]}), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_40446f2e_instance_RESULT));
assign RESULT=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_40446f2e_instance_RESULT;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_40446f2e_(GO, port_3bf115d5_, RESULT);
input		GO;
input	[15:0]	port_3bf115d5_;
output	[15:0]	RESULT;
wire signed	[15:0]	greaterThan_a_signed;
wire		greaterThan;
wire signed	[15:0]	greaterThan_b_signed;
wire		and_u187_u0;
wire		not_u36_u0;
wire		and_u188_u0;
wire		and_u189_u0;
wire		and_u190_u0;
wire	[15:0]	mux_u13;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_3bf115d5_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign and_u187_u0=GO&greaterThan;
assign not_u36_u0=~greaterThan;
assign and_u188_u0=GO&not_u36_u0;
assign and_u189_u0=and_u188_u0&GO;
assign and_u190_u0=and_u187_u0&GO;
assign mux_u13=(and_u189_u0)?port_3bf115d5_:16'h0;
assign RESULT=mux_u13;
endmodule



module LL1_H_iunzipFilter2D_endianswapper_5a2ed3eb_(endianswapper_5a2ed3eb_in, endianswapper_5a2ed3eb_out);
input	[15:0]	endianswapper_5a2ed3eb_in;
output	[15:0]	endianswapper_5a2ed3eb_out;
assign endianswapper_5a2ed3eb_out=endianswapper_5a2ed3eb_in;
endmodule



module LL1_H_iunzipFilter2D_endianswapper_28a45f1b_(endianswapper_28a45f1b_in, endianswapper_28a45f1b_out);
input	[15:0]	endianswapper_28a45f1b_in;
output	[15:0]	endianswapper_28a45f1b_out;
assign endianswapper_28a45f1b_out=endianswapper_28a45f1b_in;
endmodule



module LL1_H_iunzipFilter2D_stateVar_midPtr(bus_3400e46f_, bus_7a165d5a_, bus_538c7874_, bus_28a8a022_, bus_7badf2be_, bus_101c6579_, bus_5c59d90c_, bus_1161e5a4_, bus_64256bdd_, bus_330204f5_, bus_38b992ab_, bus_32076783_, bus_5a6e6bb4_, bus_4d247641_, bus_7ed2fb60_, bus_65180804_, bus_1be8c6a2_, bus_32f3848c_, bus_5c9b2897_, bus_123ed54b_, bus_4f392724_, bus_28004d89_, bus_7f3f31fb_, bus_1ba98a29_, bus_2d59721d_, bus_347ba71a_, bus_001a5c18_, bus_2eaf6154_, bus_32667a0e_, bus_0a10ed77_, bus_1bfd9163_, bus_4d20b648_, bus_7151a5ac_, bus_4daa9a66_, bus_35aa0d29_, bus_2ecb039d_, bus_5730d21a_, bus_48668b00_, bus_1910cc4e_, bus_6613fb43_, bus_3ae651af_, bus_53fb8955_, bus_2235ebf1_, bus_5a82cd0e_, bus_5ad36c45_);
input		bus_3400e46f_;
input		bus_7a165d5a_;
input		bus_538c7874_;
input	[15:0]	bus_28a8a022_;
input		bus_7badf2be_;
input	[15:0]	bus_101c6579_;
input		bus_5c59d90c_;
input	[15:0]	bus_1161e5a4_;
input		bus_64256bdd_;
input	[15:0]	bus_330204f5_;
input		bus_38b992ab_;
input	[15:0]	bus_32076783_;
input		bus_5a6e6bb4_;
input	[15:0]	bus_4d247641_;
input		bus_7ed2fb60_;
input	[15:0]	bus_65180804_;
input		bus_1be8c6a2_;
input	[15:0]	bus_32f3848c_;
input		bus_5c9b2897_;
input	[15:0]	bus_123ed54b_;
input		bus_4f392724_;
input	[15:0]	bus_28004d89_;
input		bus_7f3f31fb_;
input	[15:0]	bus_1ba98a29_;
input		bus_2d59721d_;
input	[15:0]	bus_347ba71a_;
input		bus_001a5c18_;
input	[15:0]	bus_2eaf6154_;
input		bus_32667a0e_;
input	[15:0]	bus_0a10ed77_;
input		bus_1bfd9163_;
input	[15:0]	bus_4d20b648_;
input		bus_7151a5ac_;
input	[15:0]	bus_4daa9a66_;
input		bus_35aa0d29_;
input	[15:0]	bus_2ecb039d_;
input		bus_5730d21a_;
input	[15:0]	bus_48668b00_;
input		bus_1910cc4e_;
input	[15:0]	bus_6613fb43_;
input		bus_3ae651af_;
input	[15:0]	bus_53fb8955_;
input		bus_2235ebf1_;
input	[15:0]	bus_5a82cd0e_;
output	[15:0]	bus_5ad36c45_;
wire	[15:0]	mux_2488d93d_u0;
wire	[15:0]	endianswapper_5a2ed3eb_out;
reg	[15:0]	stateVar_midPtr_u0=16'h0;
wire		or_71f22ffb_u0;
wire	[15:0]	endianswapper_28a45f1b_out;
assign bus_5ad36c45_=endianswapper_28a45f1b_out;
assign mux_2488d93d_u0=({16{bus_538c7874_}}&bus_28a8a022_)|({16{bus_7badf2be_}}&bus_101c6579_)|({16{bus_5c59d90c_}}&16'h0)|({16{bus_64256bdd_}}&bus_330204f5_)|({16{bus_38b992ab_}}&bus_32076783_)|({16{bus_5a6e6bb4_}}&bus_4d247641_)|({16{bus_7ed2fb60_}}&bus_65180804_)|({16{bus_1be8c6a2_}}&bus_32f3848c_)|({16{bus_5c9b2897_}}&bus_123ed54b_)|({16{bus_4f392724_}}&bus_28004d89_)|({16{bus_7f3f31fb_}}&bus_1ba98a29_)|({16{bus_2d59721d_}}&16'h0)|({16{bus_001a5c18_}}&16'h0)|({16{bus_32667a0e_}}&16'h0)|({16{bus_1bfd9163_}}&16'h0)|({16{bus_7151a5ac_}}&bus_4daa9a66_)|({16{bus_35aa0d29_}}&bus_2ecb039d_)|({16{bus_5730d21a_}}&bus_48668b00_)|({16{bus_1910cc4e_}}&bus_6613fb43_)|({16{bus_3ae651af_}}&16'h0)|({16{bus_2235ebf1_}}&16'h0);
LL1_H_iunzipFilter2D_endianswapper_5a2ed3eb_ LL1_H_iunzipFilter2D_endianswapper_5a2ed3eb__1(.endianswapper_5a2ed3eb_in(mux_2488d93d_u0), 
  .endianswapper_5a2ed3eb_out(endianswapper_5a2ed3eb_out));
always @(posedge bus_3400e46f_ or posedge bus_7a165d5a_)
begin
if (bus_7a165d5a_)
stateVar_midPtr_u0<=16'h0;
else if (or_71f22ffb_u0)
stateVar_midPtr_u0<=endianswapper_5a2ed3eb_out;
end
assign or_71f22ffb_u0=bus_538c7874_|bus_7badf2be_|bus_5c59d90c_|bus_64256bdd_|bus_38b992ab_|bus_5a6e6bb4_|bus_7ed2fb60_|bus_1be8c6a2_|bus_5c9b2897_|bus_4f392724_|bus_7f3f31fb_|bus_2d59721d_|bus_001a5c18_|bus_32667a0e_|bus_1bfd9163_|bus_7151a5ac_|bus_35aa0d29_|bus_5730d21a_|bus_1910cc4e_|bus_3ae651af_|bus_2235ebf1_;
LL1_H_iunzipFilter2D_endianswapper_28a45f1b_ LL1_H_iunzipFilter2D_endianswapper_28a45f1b__1(.endianswapper_28a45f1b_in(stateVar_midPtr_u0), 
  .endianswapper_28a45f1b_out(endianswapper_28a45f1b_out));
endmodule



module LL1_H_iunzipFilter2D_simplememoryreferee_50b1249c_(bus_3d99ccb2_, bus_4561f8d0_, bus_699bc1b7_, bus_5bec3b7f_, bus_66b004a1_, bus_3c867f89_, bus_188ca39b_, bus_315688d8_, bus_7d411a66_, bus_2da7af10_, bus_624df4b1_, bus_3fffd7cb_, bus_77051f23_, bus_3681a366_);
input		bus_3d99ccb2_;
input		bus_4561f8d0_;
input		bus_699bc1b7_;
input	[15:0]	bus_5bec3b7f_;
input		bus_66b004a1_;
input	[15:0]	bus_3c867f89_;
input	[31:0]	bus_188ca39b_;
input	[2:0]	bus_315688d8_;
output	[15:0]	bus_7d411a66_;
output	[31:0]	bus_2da7af10_;
output		bus_624df4b1_;
output		bus_3fffd7cb_;
output	[2:0]	bus_77051f23_;
output		bus_3681a366_;
assign bus_7d411a66_=bus_3c867f89_;
assign bus_2da7af10_=bus_188ca39b_;
assign bus_624df4b1_=bus_66b004a1_;
assign bus_3fffd7cb_=bus_66b004a1_;
assign bus_77051f23_=3'h1;
assign bus_3681a366_=bus_699bc1b7_;
endmodule



module LL1_H_iunzipFilter2D_midLeft1(CLK, RESET, GO, port_7c96fb9c_, port_193dec0c_, port_3a87bf5f_, port_76f10329_, port_32ad3201_, port_13cf03ae_, port_718237b9_, RESULT, RESULT_u123, RESULT_u124, RESULT_u125, RESULT_u126, RESULT_u127, RESULT_u128, RESULT_u129, RESULT_u130, RESULT_u131, RESULT_u132, RESULT_u133, RESULT_u134, RESULT_u135, RESULT_u136, RESULT_u137, RESULT_u138, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_7c96fb9c_;
input	[31:0]	port_193dec0c_;
input	[15:0]	port_3a87bf5f_;
input		port_76f10329_;
input	[15:0]	port_32ad3201_;
input		port_13cf03ae_;
input	[15:0]	port_718237b9_;
output		RESULT;
output	[15:0]	RESULT_u123;
output		RESULT_u124;
output	[31:0]	RESULT_u125;
output		RESULT_u126;
output	[15:0]	RESULT_u127;
output		RESULT_u128;
output	[31:0]	RESULT_u129;
output	[2:0]	RESULT_u130;
output		RESULT_u131;
output	[31:0]	RESULT_u132;
output	[15:0]	RESULT_u133;
output	[2:0]	RESULT_u134;
output		RESULT_u135;
output	[15:0]	RESULT_u136;
output		RESULT_u137;
output	[15:0]	RESULT_u138;
output		DONE;
wire		simplePinWrite;
wire		or_u39_u0;
wire		and_u192_u0;
reg		done_cache_u12=1'h0;
wire		or_u40_u0;
wire		and_u197_u0;
reg		done_cache_u13_u0=1'h0;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_3d0b186f_instance_RESULT;
wire		and_u206_u0;
reg		reg_64d66cce_u0=1'h0;
wire		or_u41_u0;
wire	[31:0]	add;
wire	[15:0]	add_u1;
wire		simplePinWrite_u41;
wire	[15:0]	simplePinWrite_u42;
wire	[15:0]	simplePinWrite_u43;
reg		reg_2d62db4a_u0=1'h0;
reg		reg_79ae98ce_u0=1'h0;
reg		reg_67616312_u0=1'h0;
reg	[15:0]	syncEnable_u7=16'h0;
reg		reg_6c407df9_u0=1'h0;
reg		reg_2d62db4a_result_delayed_u0=1'h0;
wire		or_u42_u0;
reg	[15:0]	syncEnable_u8_u0=16'h0;
reg		reg_6c407df9_result_delayed_u0=1'h0;
assign simplePinWrite=GO&{1{GO}};
assign or_u39_u0=and_u192_u0|RESET;
assign and_u192_u0=done_cache_u12&port_13cf03ae_;
always @(posedge CLK or posedge GO or posedge or_u39_u0)
begin
if (or_u39_u0)
done_cache_u12<=1'h0;
else if (GO)
done_cache_u12<=1'h1;
else done_cache_u12<=done_cache_u12;
end
assign or_u40_u0=and_u197_u0|RESET;
assign and_u197_u0=done_cache_u13_u0&port_13cf03ae_;
always @(posedge CLK or posedge reg_6c407df9_result_delayed_u0 or posedge or_u40_u0)
begin
if (or_u40_u0)
done_cache_u13_u0<=1'h0;
else if (reg_6c407df9_result_delayed_u0)
done_cache_u13_u0<=1'h1;
else done_cache_u13_u0<=done_cache_u13_u0;
end
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_3d0b186f_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_3d0b186f_instance(.GO(reg_79ae98ce_u0), 
  .port_1f044053_(syncEnable_u8_u0), .port_7b52a31d_(port_32ad3201_), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_3d0b186f_instance_RESULT));
assign and_u206_u0=reg_64d66cce_u0&port_13cf03ae_;
always @(posedge CLK or posedge reg_2d62db4a_result_delayed_u0 or posedge or_u41_u0)
begin
if (or_u41_u0)
reg_64d66cce_u0<=1'h0;
else if (reg_2d62db4a_result_delayed_u0)
reg_64d66cce_u0<=1'h1;
else reg_64d66cce_u0<=reg_64d66cce_u0;
end
assign or_u41_u0=and_u206_u0|RESET;
assign add=port_193dec0c_+32'h1;
assign add_u1=port_3a87bf5f_+16'h1;
assign simplePinWrite_u41=reg_79ae98ce_u0&{1{reg_79ae98ce_u0}};
assign simplePinWrite_u42=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_3d0b186f_instance_RESULT&{16{reg_79ae98ce_u0}};
assign simplePinWrite_u43=16'h1&{16{1'h1}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2d62db4a_u0<=1'h0;
else reg_2d62db4a_u0<=reg_79ae98ce_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_79ae98ce_u0<=1'h0;
else reg_79ae98ce_u0<=reg_6c407df9_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_67616312_u0<=1'h0;
else reg_67616312_u0<=reg_2d62db4a_result_delayed_u0;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u7<=port_718237b9_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6c407df9_u0<=1'h0;
else reg_6c407df9_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2d62db4a_result_delayed_u0<=1'h0;
else reg_2d62db4a_result_delayed_u0<=reg_2d62db4a_u0;
end
assign or_u42_u0=GO|reg_6c407df9_result_delayed_u0;
always @(posedge CLK)
begin
if (reg_6c407df9_u0)
syncEnable_u8_u0<=port_32ad3201_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6c407df9_result_delayed_u0<=1'h0;
else reg_6c407df9_result_delayed_u0<=reg_6c407df9_u0;
end
assign RESULT=GO;
assign RESULT_u123=16'h0;
assign RESULT_u124=GO;
assign RESULT_u125=add;
assign RESULT_u126=GO;
assign RESULT_u127=add_u1;
assign RESULT_u128=or_u42_u0;
assign RESULT_u129=32'h0;
assign RESULT_u130=3'h1;
assign RESULT_u131=reg_2d62db4a_result_delayed_u0;
assign RESULT_u132=32'h0;
assign RESULT_u133=syncEnable_u7;
assign RESULT_u134=3'h1;
assign RESULT_u135=simplePinWrite;
assign RESULT_u136=simplePinWrite_u43;
assign RESULT_u137=simplePinWrite_u41;
assign RESULT_u138=simplePinWrite_u42;
assign DONE=reg_67616312_u0;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_3d0b186f_(GO, port_1f044053_, port_7b52a31d_, RESULT);
input		GO;
input	[15:0]	port_1f044053_;
input	[15:0]	port_7b52a31d_;
output	[15:0]	RESULT;
wire	[16:0]	add;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_4935f088_instance_RESULT;
assign add={port_1f044053_[15], port_1f044053_}+{port_7b52a31d_[15], port_7b52a31d_};
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_4935f088_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_4935f088_instance(.GO(GO), 
  .port_6eff38c6_({add[16], add[16:2]}), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_4935f088_instance_RESULT));
assign RESULT=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_4935f088_instance_RESULT;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_4935f088_(GO, port_6eff38c6_, RESULT);
input		GO;
input	[15:0]	port_6eff38c6_;
output	[15:0]	RESULT;
wire signed	[15:0]	greaterThan_b_signed;
wire signed	[15:0]	greaterThan_a_signed;
wire		greaterThan;
wire		and_u201_u0;
wire		and_u202_u0;
wire		not_u37_u0;
wire		and_u203_u0;
wire		and_u204_u0;
wire	[15:0]	mux_u14;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_6eff38c6_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign and_u201_u0=GO&greaterThan;
assign and_u202_u0=GO&not_u37_u0;
assign not_u37_u0=~greaterThan;
assign and_u203_u0=and_u202_u0&GO;
assign and_u204_u0=and_u201_u0&GO;
assign mux_u14=(and_u204_u0)?16'h0:port_6eff38c6_;
assign RESULT=mux_u14;
endmodule



module LL1_H_iunzipFilter2D_Kicker_6(CLK, RESET, bus_4ae3b466_);
input		CLK;
input		RESET;
output		bus_4ae3b466_;
wire		bus_647f33a2_;
wire		bus_12d8f98f_;
reg		kicker_1=1'h0;
wire		bus_468bf43e_;
wire		bus_262977bf_;
reg		kicker_res=1'h0;
reg		kicker_2=1'h0;
assign bus_647f33a2_=~kicker_2;
assign bus_12d8f98f_=kicker_1&bus_468bf43e_&bus_647f33a2_;
always @(posedge CLK)
begin
kicker_1<=bus_468bf43e_;
end
assign bus_468bf43e_=~RESET;
assign bus_262977bf_=bus_468bf43e_&kicker_1;
always @(posedge CLK)
begin
kicker_res<=bus_12d8f98f_;
end
always @(posedge CLK)
begin
kicker_2<=bus_262977bf_;
end
assign bus_4ae3b466_=kicker_res;
endmodule



module LL1_H_iunzipFilter2D_donePopulateBuffer(CLK, RESET, GO, RESULT, RESULT_u139, DONE);
input		CLK;
input		RESET;
input		GO;
output		RESULT;
output	[15:0]	RESULT_u139;
output		DONE;
reg		reg_4beb7221_u0=1'h0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4beb7221_u0<=1'h0;
else reg_4beb7221_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u139=16'h0;
assign DONE=reg_4beb7221_u0;
endmodule



module LL1_H_iunzipFilter2D_endianswapper_2ae2ff75_(endianswapper_2ae2ff75_in, endianswapper_2ae2ff75_out);
input	[2:0]	endianswapper_2ae2ff75_in;
output	[2:0]	endianswapper_2ae2ff75_out;
assign endianswapper_2ae2ff75_out=endianswapper_2ae2ff75_in;
endmodule



module LL1_H_iunzipFilter2D_endianswapper_751a48a3_(endianswapper_751a48a3_in, endianswapper_751a48a3_out);
input	[2:0]	endianswapper_751a48a3_in;
output	[2:0]	endianswapper_751a48a3_out;
assign endianswapper_751a48a3_out=endianswapper_751a48a3_in;
endmodule



module LL1_H_iunzipFilter2D_stateVar_fsmState_LL1_H_iunzipFilter2D(bus_3aa33e9e_, bus_0f971a50_, bus_760e0512_, bus_628847e6_, bus_60d84d20_);
input		bus_3aa33e9e_;
input		bus_0f971a50_;
input		bus_760e0512_;
input	[2:0]	bus_628847e6_;
output	[2:0]	bus_60d84d20_;
wire	[2:0]	endianswapper_2ae2ff75_out;
reg	[2:0]	stateVar_fsmState_LL1_H_iunzipFilter2D_u0=3'h0;
wire	[2:0]	endianswapper_751a48a3_out;
LL1_H_iunzipFilter2D_endianswapper_2ae2ff75_ LL1_H_iunzipFilter2D_endianswapper_2ae2ff75__1(.endianswapper_2ae2ff75_in(stateVar_fsmState_LL1_H_iunzipFilter2D_u0), 
  .endianswapper_2ae2ff75_out(endianswapper_2ae2ff75_out));
always @(posedge bus_3aa33e9e_ or posedge bus_0f971a50_)
begin
if (bus_0f971a50_)
stateVar_fsmState_LL1_H_iunzipFilter2D_u0<=3'h0;
else if (bus_760e0512_)
stateVar_fsmState_LL1_H_iunzipFilter2D_u0<=endianswapper_751a48a3_out;
end
LL1_H_iunzipFilter2D_endianswapper_751a48a3_ LL1_H_iunzipFilter2D_endianswapper_751a48a3__1(.endianswapper_751a48a3_in(bus_628847e6_), 
  .endianswapper_751a48a3_out(endianswapper_751a48a3_out));
assign bus_60d84d20_=endianswapper_2ae2ff75_out;
endmodule



module LL1_H_iunzipFilter2D_bottomRightNoConsume1(CLK, RESET, GO, port_31e3635b_, port_43d1b2b6_, port_4d9c680b_, RESULT, RESULT_u140, RESULT_u141, RESULT_u142, RESULT_u143, RESULT_u144, RESULT_u145, RESULT_u146, RESULT_u147, RESULT_u148, RESULT_u149, RESULT_u150, RESULT_u151, RESULT_u152, RESULT_u153, RESULT_u154, DONE);
input		CLK;
input		RESET;
input		GO;
input		port_31e3635b_;
input		port_43d1b2b6_;
input	[15:0]	port_4d9c680b_;
output		RESULT;
output	[15:0]	RESULT_u140;
output		RESULT_u141;
output	[15:0]	RESULT_u142;
output		RESULT_u143;
output	[15:0]	RESULT_u144;
output		RESULT_u145;
output	[31:0]	RESULT_u146;
output		RESULT_u147;
output		RESULT_u148;
output		RESULT_u149;
output	[31:0]	RESULT_u150;
output	[2:0]	RESULT_u151;
output	[15:0]	RESULT_u152;
output		RESULT_u153;
output	[15:0]	RESULT_u154;
output		DONE;
wire		or_u43_u0;
wire		and_u209_u0;
reg		done_cache_u14=1'h0;
reg		done_cache_u15_u0=1'h0;
wire		or_u44_u0;
wire		and_u214_u0;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_01f7d127_instance_RESULT;
wire		not_u39;
wire	[15:0]	simplePinWrite;
wire	[15:0]	simplePinWrite_u44;
wire		simplePinWrite_u45;
reg		reg_093e282b_u0=1'h0;
reg		reg_093e282b_result_delayed_u0=1'h0;
reg	[15:0]	syncEnable_u9=16'h0;
reg		reg_17bd3836_u0=1'h0;
wire		or_u45_u0;
reg		reg_118cfc23_u0=1'h0;
reg		reg_797367b9_u0=1'h0;
assign or_u43_u0=and_u209_u0|RESET;
assign and_u209_u0=done_cache_u14&port_43d1b2b6_;
always @(posedge CLK or posedge GO or posedge or_u43_u0)
begin
if (or_u43_u0)
done_cache_u14<=1'h0;
else if (GO)
done_cache_u14<=1'h1;
else done_cache_u14<=done_cache_u14;
end
always @(posedge CLK or posedge reg_118cfc23_u0 or posedge or_u44_u0)
begin
if (or_u44_u0)
done_cache_u15_u0<=1'h0;
else if (reg_118cfc23_u0)
done_cache_u15_u0<=1'h1;
else done_cache_u15_u0<=done_cache_u15_u0;
end
assign or_u44_u0=and_u214_u0|RESET;
assign and_u214_u0=done_cache_u15_u0&port_43d1b2b6_;
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_01f7d127_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_01f7d127_instance(.GO(reg_17bd3836_u0), 
  .port_1a3748a9_(port_4d9c680b_), .port_18798b8f_(syncEnable_u9), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_01f7d127_instance_RESULT));
assign not_u39=!port_31e3635b_;
assign simplePinWrite=16'h1&{16{1'h1}};
assign simplePinWrite_u44=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_01f7d127_instance_RESULT&{16{reg_17bd3836_u0}};
assign simplePinWrite_u45=reg_17bd3836_u0&{1{reg_17bd3836_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_093e282b_u0<=1'h0;
else reg_093e282b_u0<=reg_17bd3836_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_093e282b_result_delayed_u0<=1'h0;
else reg_093e282b_result_delayed_u0<=reg_093e282b_u0;
end
always @(posedge CLK)
begin
if (reg_797367b9_u0)
syncEnable_u9<=port_4d9c680b_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_17bd3836_u0<=1'h0;
else reg_17bd3836_u0<=reg_118cfc23_u0;
end
assign or_u45_u0=GO|reg_118cfc23_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_118cfc23_u0<=1'h0;
else reg_118cfc23_u0<=reg_797367b9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_797367b9_u0<=1'h0;
else reg_797367b9_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u140=16'h0;
assign RESULT_u141=GO;
assign RESULT_u142=16'h0;
assign RESULT_u143=GO;
assign RESULT_u144=16'h0;
assign RESULT_u145=GO;
assign RESULT_u146=32'h0;
assign RESULT_u147=GO;
assign RESULT_u148=not_u39;
assign RESULT_u149=or_u45_u0;
assign RESULT_u150=32'h0;
assign RESULT_u151=3'h1;
assign RESULT_u152=simplePinWrite;
assign RESULT_u153=simplePinWrite_u45;
assign RESULT_u154=simplePinWrite_u44;
assign DONE=reg_093e282b_result_delayed_u0;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_01f7d127_(GO, port_1a3748a9_, port_18798b8f_, RESULT);
input		GO;
input	[15:0]	port_1a3748a9_;
input	[15:0]	port_18798b8f_;
output	[15:0]	RESULT;
wire	[16:0]	add;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_77e7c4ff_instance_RESULT;
assign add={port_18798b8f_[15], port_18798b8f_}+{port_1a3748a9_[15], port_1a3748a9_};
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_77e7c4ff_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_77e7c4ff_instance(.GO(GO), 
  .port_063a73f3_({add[16], add[16:2]}), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_77e7c4ff_instance_RESULT));
assign RESULT=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_77e7c4ff_instance_RESULT;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_77e7c4ff_(GO, port_063a73f3_, RESULT);
input		GO;
input	[15:0]	port_063a73f3_;
output	[15:0]	RESULT;
wire		greaterThan;
wire signed	[15:0]	greaterThan_b_signed;
wire signed	[15:0]	greaterThan_a_signed;
wire		and_u218_u0;
wire		and_u219_u0;
wire		not_u38_u0;
wire	[15:0]	mux_u15;
wire		and_u220_u0;
wire		and_u221_u0;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_063a73f3_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign and_u218_u0=GO&greaterThan;
assign and_u219_u0=GO&not_u38_u0;
assign not_u38_u0=~greaterThan;
assign mux_u15=(and_u221_u0)?16'h0:port_063a73f3_;
assign and_u220_u0=and_u219_u0&GO;
assign and_u221_u0=and_u218_u0&GO;
assign RESULT=mux_u15;
endmodule



module LL1_H_iunzipFilter2D_stateVar_isEven(bus_16c94a5f_, bus_06dd97a7_, bus_23cf6553_, bus_1582983e_, bus_193ba992_, bus_250aabcd_, bus_1503fca4_, bus_052f1bad_, bus_5b66ba18_, bus_0fdbb770_, bus_64dea1fa_, bus_652c6729_, bus_4d350cfd_, bus_0dca5a75_, bus_1946dfc4_, bus_06915c78_, bus_15ebb497_);
input		bus_16c94a5f_;
input		bus_06dd97a7_;
input		bus_23cf6553_;
input		bus_1582983e_;
input		bus_193ba992_;
input		bus_250aabcd_;
input		bus_1503fca4_;
input		bus_052f1bad_;
input		bus_5b66ba18_;
input		bus_0fdbb770_;
input		bus_64dea1fa_;
input		bus_652c6729_;
input		bus_4d350cfd_;
input		bus_0dca5a75_;
input		bus_1946dfc4_;
input		bus_06915c78_;
output		bus_15ebb497_;
wire		mux_5ccbbeed_u0;
wire		or_5c83c9a5_u0;
reg		stateVar_isEven_u0=1'h1;
assign mux_5ccbbeed_u0=({1{bus_23cf6553_}}&bus_1582983e_)|({1{bus_193ba992_}}&bus_250aabcd_)|({1{bus_1503fca4_}}&bus_052f1bad_)|({1{bus_5b66ba18_}}&bus_0fdbb770_)|({1{bus_64dea1fa_}}&bus_652c6729_)|({1{bus_4d350cfd_}}&bus_0dca5a75_)|({1{bus_1946dfc4_}}&bus_06915c78_);
assign or_5c83c9a5_u0=bus_23cf6553_|bus_193ba992_|bus_1503fca4_|bus_5b66ba18_|bus_64dea1fa_|bus_4d350cfd_|bus_1946dfc4_;
always @(posedge bus_16c94a5f_ or posedge bus_06dd97a7_)
begin
if (bus_06dd97a7_)
stateVar_isEven_u0<=1'h1;
else if (or_5c83c9a5_u0)
stateVar_isEven_u0<=mux_5ccbbeed_u0;
end
assign bus_15ebb497_=stateVar_isEven_u0;
endmodule



module LL1_H_iunzipFilter2D_bottomLeftNoConsume2(CLK, RESET, GO, port_773c7b8d_, port_18be374b_, port_373fd3b4_, port_59b7d69f_, RESULT, RESULT_u155, RESULT_u156, RESULT_u157, RESULT_u158, RESULT_u159, RESULT_u160, RESULT_u161, RESULT_u162, RESULT_u163, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_773c7b8d_;
input	[15:0]	port_18be374b_;
input		port_373fd3b4_;
input	[15:0]	port_59b7d69f_;
output		RESULT;
output	[15:0]	RESULT_u155;
output		RESULT_u156;
output	[15:0]	RESULT_u157;
output		RESULT_u158;
output	[31:0]	RESULT_u159;
output	[2:0]	RESULT_u160;
output	[15:0]	RESULT_u161;
output		RESULT_u162;
output	[15:0]	RESULT_u163;
output		DONE;
wire		or_u46_u0;
reg		done_cache_u16=1'h0;
wire		and_u222_u0;
wire		or_u47_u0;
reg		done_cache_u17_u0=1'h0;
wire		and_u227_u0;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_6d3415e3_instance_RESULT;
wire	[15:0]	add;
wire		simplePinWrite;
wire	[15:0]	simplePinWrite_u46;
wire	[15:0]	simplePinWrite_u47;
reg		reg_2ce6f3d1_u0=1'h0;
reg		reg_51f5879e_u0=1'h0;
wire		or_u48_u0;
reg		reg_4a157363_u0=1'h0;
reg	[15:0]	syncEnable_u10=16'h0;
reg		reg_2ce6f3d1_result_delayed_u0=1'h0;
reg		reg_40d29a0a_u0=1'h0;
assign or_u46_u0=and_u222_u0|RESET;
always @(posedge CLK or posedge GO or posedge or_u46_u0)
begin
if (or_u46_u0)
done_cache_u16<=1'h0;
else if (GO)
done_cache_u16<=1'h1;
else done_cache_u16<=done_cache_u16;
end
assign and_u222_u0=done_cache_u16&port_373fd3b4_;
assign or_u47_u0=and_u227_u0|RESET;
always @(posedge CLK or posedge reg_51f5879e_u0 or posedge or_u47_u0)
begin
if (or_u47_u0)
done_cache_u17_u0<=1'h0;
else if (reg_51f5879e_u0)
done_cache_u17_u0<=1'h1;
else done_cache_u17_u0<=done_cache_u17_u0;
end
assign and_u227_u0=done_cache_u17_u0&port_373fd3b4_;
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_6d3415e3_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_6d3415e3_instance(.GO(reg_2ce6f3d1_u0), 
  .port_232c036f_(port_59b7d69f_), .port_6b27401f_(syncEnable_u10), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_6d3415e3_instance_RESULT));
assign add=port_18be374b_+16'h1;
assign simplePinWrite=reg_2ce6f3d1_u0&{1{reg_2ce6f3d1_u0}};
assign simplePinWrite_u46=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_6d3415e3_instance_RESULT&{16{reg_2ce6f3d1_u0}};
assign simplePinWrite_u47=16'h1&{16{1'h1}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2ce6f3d1_u0<=1'h0;
else reg_2ce6f3d1_u0<=reg_51f5879e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_51f5879e_u0<=1'h0;
else reg_51f5879e_u0<=reg_40d29a0a_u0;
end
assign or_u48_u0=GO|reg_51f5879e_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4a157363_u0<=1'h0;
else reg_4a157363_u0<=reg_2ce6f3d1_result_delayed_u0;
end
always @(posedge CLK)
begin
if (reg_40d29a0a_u0)
syncEnable_u10<=port_59b7d69f_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2ce6f3d1_result_delayed_u0<=1'h0;
else reg_2ce6f3d1_result_delayed_u0<=reg_2ce6f3d1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_40d29a0a_u0<=1'h0;
else reg_40d29a0a_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u155=16'h0;
assign RESULT_u156=GO;
assign RESULT_u157=add;
assign RESULT_u158=or_u48_u0;
assign RESULT_u159=32'h0;
assign RESULT_u160=3'h1;
assign RESULT_u161=simplePinWrite_u47;
assign RESULT_u162=simplePinWrite;
assign RESULT_u163=simplePinWrite_u46;
assign DONE=reg_4a157363_u0;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_6d3415e3_(GO, port_232c036f_, port_6b27401f_, RESULT);
input		GO;
input	[15:0]	port_232c036f_;
input	[15:0]	port_6b27401f_;
output	[15:0]	RESULT;
wire	[15:0]	subtract;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_0979a93a_instance_RESULT;
assign subtract=port_6b27401f_-port_232c036f_;
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_0979a93a_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_0979a93a_instance(.GO(GO), 
  .port_53326142_({subtract[15], subtract[15:1]}), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_0979a93a_instance_RESULT));
assign RESULT=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_0979a93a_instance_RESULT;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_0979a93a_(GO, port_53326142_, RESULT);
input		GO;
input	[15:0]	port_53326142_;
output	[15:0]	RESULT;
wire signed	[15:0]	greaterThan_b_signed;
wire signed	[15:0]	greaterThan_a_signed;
wire		greaterThan;
wire		not_u40_u0;
wire		and_u231_u0;
wire		and_u232_u0;
wire	[15:0]	mux_u16;
wire		and_u233_u0;
wire		and_u234_u0;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_53326142_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign not_u40_u0=~greaterThan;
assign and_u231_u0=GO&greaterThan;
assign and_u232_u0=GO&not_u40_u0;
assign mux_u16=(and_u233_u0)?16'h0:port_53326142_;
assign and_u233_u0=and_u231_u0&GO;
assign and_u234_u0=and_u232_u0&GO;
assign RESULT=mux_u16;
endmodule



module LL1_H_iunzipFilter2D_topLeft(CLK, RESET, GO, port_5221a8c5_, port_2026972c_, port_6d155da5_, port_792b0e97_, port_20f4db23_, port_50f97c55_, port_6e419463_, RESULT, RESULT_u164, RESULT_u165, RESULT_u166, RESULT_u167, RESULT_u168, RESULT_u169, RESULT_u170, RESULT_u171, RESULT_u172, RESULT_u173, RESULT_u174, RESULT_u175, RESULT_u176, RESULT_u177, RESULT_u178, RESULT_u179, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_5221a8c5_;
input	[31:0]	port_2026972c_;
input	[15:0]	port_6d155da5_;
input		port_792b0e97_;
input	[15:0]	port_20f4db23_;
input		port_50f97c55_;
input	[15:0]	port_6e419463_;
output		RESULT;
output	[15:0]	RESULT_u164;
output		RESULT_u165;
output	[31:0]	RESULT_u166;
output		RESULT_u167;
output	[15:0]	RESULT_u168;
output		RESULT_u169;
output	[31:0]	RESULT_u170;
output	[2:0]	RESULT_u171;
output		RESULT_u172;
output	[31:0]	RESULT_u173;
output	[15:0]	RESULT_u174;
output	[2:0]	RESULT_u175;
output		RESULT_u176;
output	[15:0]	RESULT_u177;
output		RESULT_u178;
output	[15:0]	RESULT_u179;
output		DONE;
wire		simplePinWrite;
wire		and_u236_u0;
wire		or_u49_u0;
reg		done_cache_u18=1'h0;
wire		or_u50_u0;
wire		and_u239_u0;
reg		done_cache_u19_u0=1'h0;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_2a5573fa_instance_RESULT;
wire	[31:0]	add;
reg		reg_761d558d_u0=1'h0;
wire		or_u51_u0;
wire		and_u247_u0;
wire	[15:0]	add_u2;
wire	[31:0]	add_u3;
wire	[15:0]	simplePinWrite_u48;
wire	[15:0]	simplePinWrite_u49;
wire		simplePinWrite_u50;
reg		reg_5bd2a0f6_u0=1'h0;
reg	[15:0]	syncEnable_u11=16'h0;
reg		reg_5523b66a_u0=1'h0;
reg		reg_002ee37c_u0=1'h0;
reg	[31:0]	syncEnable_u12_u0=32'h0;
reg		reg_0ed6c6af_u0=1'h0;
reg	[15:0]	syncEnable_u13_u0=16'h0;
reg		reg_002ee37c_result_delayed_u0=1'h0;
reg		reg_5bd2a0f6_result_delayed_u0=1'h0;
wire	[31:0]	mux_u18;
wire		or_u52_u0;
assign simplePinWrite=GO&{1{GO}};
assign and_u236_u0=done_cache_u18&port_50f97c55_;
assign or_u49_u0=and_u236_u0|RESET;
always @(posedge CLK or posedge GO or posedge or_u49_u0)
begin
if (or_u49_u0)
done_cache_u18<=1'h0;
else if (GO)
done_cache_u18<=1'h1;
else done_cache_u18<=done_cache_u18;
end
assign or_u50_u0=and_u239_u0|RESET;
assign and_u239_u0=done_cache_u19_u0&port_50f97c55_;
always @(posedge CLK or posedge reg_5bd2a0f6_result_delayed_u0 or posedge or_u50_u0)
begin
if (or_u50_u0)
done_cache_u19_u0<=1'h0;
else if (reg_5bd2a0f6_result_delayed_u0)
done_cache_u19_u0<=1'h1;
else done_cache_u19_u0<=done_cache_u19_u0;
end
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_2a5573fa_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_2a5573fa_instance(.GO(reg_002ee37c_u0), 
  .port_1d9b49c5_(syncEnable_u11), .port_58f76ace_(port_20f4db23_), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_2a5573fa_instance_RESULT));
assign add=port_2026972c_+32'h0;
always @(posedge CLK or posedge reg_0ed6c6af_u0 or posedge or_u51_u0)
begin
if (or_u51_u0)
reg_761d558d_u0<=1'h0;
else if (reg_0ed6c6af_u0)
reg_761d558d_u0<=1'h1;
else reg_761d558d_u0<=reg_761d558d_u0;
end
assign or_u51_u0=and_u247_u0|RESET;
assign and_u247_u0=reg_761d558d_u0&port_50f97c55_;
assign add_u2=port_6d155da5_+16'h1;
assign add_u3=port_2026972c_+32'h1;
assign simplePinWrite_u48=16'h1&{16{1'h1}};
assign simplePinWrite_u49=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_2a5573fa_instance_RESULT&{16{reg_002ee37c_u0}};
assign simplePinWrite_u50=reg_002ee37c_u0&{1{reg_002ee37c_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5bd2a0f6_u0<=1'h0;
else reg_5bd2a0f6_u0<=GO;
end
always @(posedge CLK)
begin
if (reg_5bd2a0f6_u0)
syncEnable_u11<=port_20f4db23_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5523b66a_u0<=1'h0;
else reg_5523b66a_u0<=reg_0ed6c6af_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_002ee37c_u0<=1'h0;
else reg_002ee37c_u0<=reg_5bd2a0f6_result_delayed_u0;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u12_u0<=add;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0ed6c6af_u0<=1'h0;
else reg_0ed6c6af_u0<=reg_002ee37c_result_delayed_u0;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u13_u0<=port_6e419463_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_002ee37c_result_delayed_u0<=1'h0;
else reg_002ee37c_result_delayed_u0<=reg_002ee37c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5bd2a0f6_result_delayed_u0<=1'h0;
else reg_5bd2a0f6_result_delayed_u0<=reg_5bd2a0f6_u0;
end
assign mux_u18=({32{reg_0ed6c6af_u0}}&syncEnable_u12_u0)|({32{GO}}&32'h0)|({32{reg_5bd2a0f6_result_delayed_u0}}&32'h0);
assign or_u52_u0=GO|reg_5bd2a0f6_result_delayed_u0;
assign RESULT=GO;
assign RESULT_u164=16'h0;
assign RESULT_u165=GO;
assign RESULT_u166=add_u3;
assign RESULT_u167=GO;
assign RESULT_u168=add_u2;
assign RESULT_u169=or_u52_u0;
assign RESULT_u170=mux_u18;
assign RESULT_u171=3'h1;
assign RESULT_u172=reg_0ed6c6af_u0;
assign RESULT_u173=mux_u18;
assign RESULT_u174=syncEnable_u13_u0;
assign RESULT_u175=3'h1;
assign RESULT_u176=simplePinWrite;
assign RESULT_u177=simplePinWrite_u48;
assign RESULT_u178=simplePinWrite_u50;
assign RESULT_u179=simplePinWrite_u49;
assign DONE=reg_5523b66a_u0;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_2a5573fa_(GO, port_1d9b49c5_, port_58f76ace_, RESULT);
input		GO;
input	[15:0]	port_1d9b49c5_;
input	[15:0]	port_58f76ace_;
output	[15:0]	RESULT;
wire	[16:0]	add;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_3f772e5c_instance_RESULT;
assign add={port_1d9b49c5_[15], port_1d9b49c5_}+{port_58f76ace_[15], port_58f76ace_};
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_3f772e5c_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_3f772e5c_instance(.GO(GO), 
  .port_132bd03d_({add[16], add[16:2]}), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_3f772e5c_instance_RESULT));
assign RESULT=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_3f772e5c_instance_RESULT;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_3f772e5c_(GO, port_132bd03d_, RESULT);
input		GO;
input	[15:0]	port_132bd03d_;
output	[15:0]	RESULT;
wire signed	[15:0]	greaterThan_b_signed;
wire signed	[15:0]	greaterThan_a_signed;
wire		greaterThan;
wire		not_u41_u0;
wire		and_u243_u0;
wire		and_u244_u0;
wire		and_u245_u0;
wire	[15:0]	mux_u17;
wire		and_u246_u0;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_132bd03d_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign not_u41_u0=~greaterThan;
assign and_u243_u0=GO&greaterThan;
assign and_u244_u0=GO&not_u41_u0;
assign and_u245_u0=and_u243_u0&GO;
assign mux_u17=(and_u245_u0)?16'h0:port_132bd03d_;
assign and_u246_u0=and_u244_u0&GO;
assign RESULT=mux_u17;
endmodule



module LL1_H_iunzipFilter2D_topRight(CLK, RESET, GO, port_21a33c82_, port_1f205dca_, port_468f8c2d_, port_05847a01_, port_0a351222_, port_19cb6266_, RESULT, RESULT_u180, RESULT_u181, RESULT_u182, RESULT_u183, RESULT_u184, RESULT_u185, RESULT_u186, RESULT_u187, RESULT_u188, RESULT_u189, RESULT_u190, RESULT_u191, RESULT_u192, RESULT_u193, RESULT_u194, RESULT_u195, RESULT_u196, RESULT_u197, RESULT_u198, RESULT_u199, DONE);
input		CLK;
input		RESET;
input		GO;
input	[31:0]	port_21a33c82_;
input		port_1f205dca_;
input		port_468f8c2d_;
input	[15:0]	port_05847a01_;
input		port_0a351222_;
input	[15:0]	port_19cb6266_;
output		RESULT;
output	[31:0]	RESULT_u180;
output		RESULT_u181;
output	[15:0]	RESULT_u182;
output		RESULT_u183;
output	[15:0]	RESULT_u184;
output		RESULT_u185;
output	[15:0]	RESULT_u186;
output		RESULT_u187;
output		RESULT_u188;
output		RESULT_u189;
output	[31:0]	RESULT_u190;
output	[2:0]	RESULT_u191;
output		RESULT_u192;
output	[31:0]	RESULT_u193;
output	[15:0]	RESULT_u194;
output	[2:0]	RESULT_u195;
output		RESULT_u196;
output	[15:0]	RESULT_u197;
output		RESULT_u198;
output	[15:0]	RESULT_u199;
output		DONE;
wire		simplePinWrite;
wire		and_u250_u0;
wire		or_u53_u0;
reg		done_cache_u20=1'h0;
wire		or_u54_u0;
wire		and_u254_u0;
reg		done_cache_u21_u0=1'h0;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_2f405190_instance_RESULT;
reg		reg_4a2406c5_u0=1'h0;
wire		and_u263_u0;
wire		or_u55_u0;
wire	[31:0]	add;
wire		not_u43;
wire	[15:0]	simplePinWrite_u51;
wire		simplePinWrite_u52;
wire	[15:0]	simplePinWrite_u53;
wire		or_u56_u0;
reg		reg_4dfa39e0_u0=1'h0;
reg	[15:0]	syncEnable_u14=16'h0;
reg		reg_317ea2fa_u0=1'h0;
reg		reg_65a68b72_u0=1'h0;
reg		reg_317ea2fa_result_delayed_u0=1'h0;
reg		reg_2a751396_u0=1'h0;
reg	[15:0]	syncEnable_u15_u0=16'h0;
reg		reg_4dfa39e0_result_delayed_u0=1'h0;
assign simplePinWrite=GO&{1{GO}};
assign and_u250_u0=done_cache_u20&port_0a351222_;
assign or_u53_u0=and_u250_u0|RESET;
always @(posedge CLK or posedge GO or posedge or_u53_u0)
begin
if (or_u53_u0)
done_cache_u20<=1'h0;
else if (GO)
done_cache_u20<=1'h1;
else done_cache_u20<=done_cache_u20;
end
assign or_u54_u0=and_u254_u0|RESET;
assign and_u254_u0=done_cache_u21_u0&port_0a351222_;
always @(posedge CLK or posedge reg_4dfa39e0_u0 or posedge or_u54_u0)
begin
if (or_u54_u0)
done_cache_u21_u0<=1'h0;
else if (reg_4dfa39e0_u0)
done_cache_u21_u0<=1'h1;
else done_cache_u21_u0<=done_cache_u21_u0;
end
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_2f405190_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_2f405190_instance(.GO(reg_4dfa39e0_result_delayed_u0), 
  .port_0e9f4280_(syncEnable_u15_u0), .port_4fef298e_(port_05847a01_), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_2f405190_instance_RESULT));
always @(posedge CLK or posedge reg_317ea2fa_result_delayed_u0 or posedge or_u55_u0)
begin
if (or_u55_u0)
reg_4a2406c5_u0<=1'h0;
else if (reg_317ea2fa_result_delayed_u0)
reg_4a2406c5_u0<=1'h1;
else reg_4a2406c5_u0<=reg_4a2406c5_u0;
end
assign and_u263_u0=reg_4a2406c5_u0&port_0a351222_;
assign or_u55_u0=and_u263_u0|RESET;
assign add=port_21a33c82_+32'h1;
assign not_u43=!port_1f205dca_;
assign simplePinWrite_u51=16'h1&{16{1'h1}};
assign simplePinWrite_u52=reg_4dfa39e0_result_delayed_u0&{1{reg_4dfa39e0_result_delayed_u0}};
assign simplePinWrite_u53=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_2f405190_instance_RESULT&{16{reg_4dfa39e0_result_delayed_u0}};
assign or_u56_u0=GO|reg_4dfa39e0_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4dfa39e0_u0<=1'h0;
else reg_4dfa39e0_u0<=reg_2a751396_u0;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u14<=port_19cb6266_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_317ea2fa_u0<=1'h0;
else reg_317ea2fa_u0<=reg_4dfa39e0_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_65a68b72_u0<=1'h0;
else reg_65a68b72_u0<=reg_317ea2fa_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_317ea2fa_result_delayed_u0<=1'h0;
else reg_317ea2fa_result_delayed_u0<=reg_317ea2fa_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2a751396_u0<=1'h0;
else reg_2a751396_u0<=GO;
end
always @(posedge CLK)
begin
if (reg_2a751396_u0)
syncEnable_u15_u0<=port_05847a01_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4dfa39e0_result_delayed_u0<=1'h0;
else reg_4dfa39e0_result_delayed_u0<=reg_4dfa39e0_u0;
end
assign RESULT=GO;
assign RESULT_u180=add;
assign RESULT_u181=GO;
assign RESULT_u182=16'h0;
assign RESULT_u183=GO;
assign RESULT_u184=16'h0;
assign RESULT_u185=GO;
assign RESULT_u186=16'h1;
assign RESULT_u187=GO;
assign RESULT_u188=not_u43;
assign RESULT_u189=or_u56_u0;
assign RESULT_u190=32'h0;
assign RESULT_u191=3'h1;
assign RESULT_u192=reg_317ea2fa_result_delayed_u0;
assign RESULT_u193=32'h0;
assign RESULT_u194=syncEnable_u14;
assign RESULT_u195=3'h1;
assign RESULT_u196=simplePinWrite;
assign RESULT_u197=simplePinWrite_u51;
assign RESULT_u198=simplePinWrite_u52;
assign RESULT_u199=simplePinWrite_u53;
assign DONE=reg_65a68b72_u0;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_2f405190_(GO, port_0e9f4280_, port_4fef298e_, RESULT);
input		GO;
input	[15:0]	port_0e9f4280_;
input	[15:0]	port_4fef298e_;
output	[15:0]	RESULT;
wire	[16:0]	add;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_4bf36956_instance_RESULT;
assign add={port_0e9f4280_[15], port_0e9f4280_}+{port_4fef298e_[15], port_4fef298e_};
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_4bf36956_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_4bf36956_instance(.GO(GO), 
  .port_7dce836c_({add[16], add[16:2]}), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_4bf36956_instance_RESULT));
assign RESULT=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_4bf36956_instance_RESULT;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_4bf36956_(GO, port_7dce836c_, RESULT);
input		GO;
input	[15:0]	port_7dce836c_;
output	[15:0]	RESULT;
wire signed	[15:0]	greaterThan_b_signed;
wire signed	[15:0]	greaterThan_a_signed;
wire		greaterThan;
wire		not_u42_u0;
wire		and_u258_u0;
wire		and_u259_u0;
wire		and_u260_u0;
wire	[15:0]	mux_u19;
wire		and_u261_u0;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_7dce836c_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign not_u42_u0=~greaterThan;
assign and_u258_u0=GO&greaterThan;
assign and_u259_u0=GO&not_u42_u0;
assign and_u260_u0=and_u259_u0&GO;
assign mux_u19=(and_u260_u0)?port_7dce836c_:16'h0;
assign and_u261_u0=and_u258_u0&GO;
assign RESULT=mux_u19;
endmodule



module LL1_H_iunzipFilter2D_forge_memory_515x16_1(CLK, ENA, WEA, DINA, ENB, WEB, DINB, ADDRA, ADDRB, DOUTA, DOUTB, DONEA, DONEB);
input		CLK;
input		ENA;
input		WEA;
input	[15:0]	DINA;
input		ENB;
input		WEB;
input	[15:0]	DINB;
input	[31:0]	ADDRA;
input	[31:0]	ADDRB;
output	[15:0]	DOUTA;
output	[15:0]	DOUTB;
output		DONEA;
output		DONEB;
wire		wea_0;
wire		web_0;
wire	[15:0]	pre_douta_0;
wire	[15:0]	pre_doutb_0;
wire	[1:0]	extrasa_0;
wire	[1:0]	extrasb_0;
reg	[15:0]	mux_outa;
reg	[15:0]	mux_outb;
reg	[31:0]	ADDRA_reg;
reg	[31:0]	ADDRB_reg;
reg		reb_done;
reg		wea_done;
reg		web_done;
reg		rea_done;
assign wea_0=WEA&(ADDRA[31:10]==22'h0);
assign web_0=WEB&(ADDRB[31:10]==22'h0);
always @(posedge CLK)
begin
ADDRA_reg<=ADDRA;
end
always @(pre_douta_0)
begin
mux_outa<=pre_douta_0;
end
always @(posedge CLK)
begin
ADDRB_reg<=ADDRB;
end
always @(pre_doutb_0)
begin
mux_outb<=pre_doutb_0;
end
always @(posedge CLK)
begin
wea_done<=WEA;
rea_done<=ENA;
web_done<=WEB;
reb_done<=ENB;
end
assign DONEA=wea_done|rea_done;
assign DONEB=web_done|reb_done;
assign DOUTA=mux_outa;
assign DOUTB=mux_outb;
// Memory array element: COL: 0, ROW: 0
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S18_S18#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S18_S18_instance_0(.CLKA(CLK), 
  .WEA(wea_0), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[15:0]), .DOA(pre_douta_0[15:0]), 
  .DIPA(2'b0), .DOPA(), .CLKB(CLK), .WEB(web_0), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), 
  .DIB(DINB[15:0]), .DOB(pre_doutb_0[15:0]), .DIPB(2'b0), .DOPB());
endmodule



module LL1_H_iunzipFilter2D_structuralmemory_7648df26_(CLK_u0, bus_7be93387_, bus_500680a1_, bus_14ede39e_, bus_6f816ba1_, bus_06d1faa7_, bus_2ac66d9a_, bus_4cb922b4_, bus_7077ea2b_, bus_2b14349a_, bus_6e848c4c_, bus_6da7b786_, bus_25361c61_, bus_02cec1f3_, bus_6dd7c8fd_, bus_7faecdeb_);
input		CLK_u0;
input		bus_7be93387_;
input	[31:0]	bus_500680a1_;
input	[2:0]	bus_14ede39e_;
input		bus_6f816ba1_;
input		bus_06d1faa7_;
input	[15:0]	bus_2ac66d9a_;
input	[31:0]	bus_4cb922b4_;
input	[2:0]	bus_7077ea2b_;
input		bus_2b14349a_;
input		bus_6e848c4c_;
input	[15:0]	bus_6da7b786_;
output	[15:0]	bus_25361c61_;
output		bus_02cec1f3_;
output	[15:0]	bus_6dd7c8fd_;
output		bus_7faecdeb_;
reg		logicalMem_5be7d2da_re_delay0_u0=1'h0;
reg		logicalMem_5be7d2da_we_delay0_u0=1'h0;
wire		or_3a4a9292_u0;
reg		logicalMem_5be7d2da_re_delay0_u1_u0=1'h0;
wire		or_1e1a06b8_u0;
wire		or_53b3a2c7_u0;
wire		or_7b78b34c_u0;
wire	[15:0]	bus_4f77e7fb_;
wire	[15:0]	bus_4e11bef2_;
reg		logicalMem_5be7d2da_we_delay0_u1_u0=1'h0;
always @(posedge CLK_u0 or posedge bus_7be93387_)
begin
if (bus_7be93387_)
logicalMem_5be7d2da_re_delay0_u0<=1'h0;
else logicalMem_5be7d2da_re_delay0_u0<=bus_2b14349a_;
end
always @(posedge CLK_u0 or posedge bus_7be93387_)
begin
if (bus_7be93387_)
logicalMem_5be7d2da_we_delay0_u0<=1'h0;
else logicalMem_5be7d2da_we_delay0_u0<=bus_06d1faa7_;
end
assign or_3a4a9292_u0=bus_6f816ba1_|bus_06d1faa7_;
always @(posedge CLK_u0 or posedge bus_7be93387_)
begin
if (bus_7be93387_)
logicalMem_5be7d2da_re_delay0_u1_u0<=1'h0;
else logicalMem_5be7d2da_re_delay0_u1_u0<=bus_6f816ba1_;
end
assign or_1e1a06b8_u0=logicalMem_5be7d2da_re_delay0_u0|logicalMem_5be7d2da_we_delay0_u1_u0;
assign bus_25361c61_=bus_4e11bef2_;
assign bus_02cec1f3_=or_53b3a2c7_u0;
assign bus_6dd7c8fd_=bus_4f77e7fb_;
assign bus_7faecdeb_=or_1e1a06b8_u0;
assign or_53b3a2c7_u0=logicalMem_5be7d2da_re_delay0_u1_u0|logicalMem_5be7d2da_we_delay0_u0;
assign or_7b78b34c_u0=bus_2b14349a_|bus_6e848c4c_;
LL1_H_iunzipFilter2D_forge_memory_515x16_1 LL1_H_iunzipFilter2D_forge_memory_515x16_1_instance0(.CLK(CLK_u0), 
  .ENA(or_3a4a9292_u0), .WEA(bus_06d1faa7_), .DINA(bus_2ac66d9a_), .ADDRA(bus_500680a1_), 
  .DOUTA(bus_4e11bef2_), .DONEA(), .ENB(or_7b78b34c_u0), .WEB(bus_6e848c4c_), .DINB(bus_6da7b786_), 
  .ADDRB(bus_4cb922b4_), .DOUTB(bus_4f77e7fb_), .DONEB());
always @(posedge CLK_u0 or posedge bus_7be93387_)
begin
if (bus_7be93387_)
logicalMem_5be7d2da_we_delay0_u1_u0<=1'h0;
else logicalMem_5be7d2da_we_delay0_u1_u0<=bus_6e848c4c_;
end
endmodule



module LL1_H_iunzipFilter2D_midNoConsume1(CLK, RESET, GO, port_45028bf7_, port_6e1d3735_, port_55325b56_, RESULT, RESULT_u200, RESULT_u201, RESULT_u202, RESULT_u203, RESULT_u204, RESULT_u205, RESULT_u206, RESULT_u207, RESULT_u208, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_45028bf7_;
input		port_6e1d3735_;
input	[15:0]	port_55325b56_;
output		RESULT;
output	[15:0]	RESULT_u200;
output		RESULT_u201;
output	[15:0]	RESULT_u202;
output		RESULT_u203;
output	[31:0]	RESULT_u204;
output	[2:0]	RESULT_u205;
output	[15:0]	RESULT_u206;
output		RESULT_u207;
output	[15:0]	RESULT_u208;
output		DONE;
wire		or_u57_u0;
reg		done_cache_u22=1'h0;
wire		and_u266_u0;
wire		and_u271_u0;
wire		or_u58_u0;
reg		done_cache_u23_u0=1'h0;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_258d1a6d_instance_RESULT;
wire	[15:0]	add;
wire	[15:0]	simplePinWrite;
wire	[15:0]	simplePinWrite_u54;
wire		simplePinWrite_u55;
wire		or_u59_u0;
reg		reg_55f833b9_u0=1'h0;
reg		reg_07d4b656_u0=1'h0;
reg		reg_191e8191_u0=1'h0;
reg		reg_55f833b9_result_delayed_u0=1'h0;
reg	[15:0]	syncEnable_u16=16'h0;
reg		reg_55f833b9_result_delayed_result_delayed_u0=1'h0;
assign or_u57_u0=and_u266_u0|RESET;
always @(posedge CLK or posedge GO or posedge or_u57_u0)
begin
if (or_u57_u0)
done_cache_u22<=1'h0;
else if (GO)
done_cache_u22<=1'h1;
else done_cache_u22<=done_cache_u22;
end
assign and_u266_u0=done_cache_u22&port_6e1d3735_;
assign and_u271_u0=done_cache_u23_u0&port_6e1d3735_;
assign or_u58_u0=and_u271_u0|RESET;
always @(posedge CLK or posedge reg_55f833b9_u0 or posedge or_u58_u0)
begin
if (or_u58_u0)
done_cache_u23_u0<=1'h0;
else if (reg_55f833b9_u0)
done_cache_u23_u0<=1'h1;
else done_cache_u23_u0<=done_cache_u23_u0;
end
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_258d1a6d_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_258d1a6d_instance(.GO(reg_55f833b9_result_delayed_u0), 
  .port_5de780e5_(syncEnable_u16), .port_70f22cc8_(port_55325b56_), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_258d1a6d_instance_RESULT));
assign add=port_45028bf7_+16'h1;
assign simplePinWrite=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_258d1a6d_instance_RESULT&{16{reg_55f833b9_result_delayed_u0}};
assign simplePinWrite_u54=16'h1&{16{1'h1}};
assign simplePinWrite_u55=reg_55f833b9_result_delayed_u0&{1{reg_55f833b9_result_delayed_u0}};
assign or_u59_u0=GO|reg_55f833b9_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_55f833b9_u0<=1'h0;
else reg_55f833b9_u0<=reg_07d4b656_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_07d4b656_u0<=1'h0;
else reg_07d4b656_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_191e8191_u0<=1'h0;
else reg_191e8191_u0<=reg_55f833b9_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_55f833b9_result_delayed_u0<=1'h0;
else reg_55f833b9_result_delayed_u0<=reg_55f833b9_u0;
end
always @(posedge CLK)
begin
if (reg_07d4b656_u0)
syncEnable_u16<=port_55325b56_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_55f833b9_result_delayed_result_delayed_u0<=1'h0;
else reg_55f833b9_result_delayed_result_delayed_u0<=reg_55f833b9_result_delayed_u0;
end
assign RESULT=GO;
assign RESULT_u200=16'h0;
assign RESULT_u201=GO;
assign RESULT_u202=add;
assign RESULT_u203=or_u59_u0;
assign RESULT_u204=32'h0;
assign RESULT_u205=3'h1;
assign RESULT_u206=simplePinWrite_u54;
assign RESULT_u207=simplePinWrite_u55;
assign RESULT_u208=simplePinWrite;
assign DONE=reg_191e8191_u0;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_258d1a6d_(GO, port_5de780e5_, port_70f22cc8_, RESULT);
input		GO;
input	[15:0]	port_5de780e5_;
input	[15:0]	port_70f22cc8_;
output	[15:0]	RESULT;
wire	[16:0]	add;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_070f4d12_instance_RESULT;
assign add={port_5de780e5_[15], port_5de780e5_}+{port_70f22cc8_[15], port_70f22cc8_};
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_070f4d12_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_070f4d12_instance(.GO(GO), 
  .port_5374d8fd_({add[16], add[16:2]}), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_070f4d12_instance_RESULT));
assign RESULT=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_070f4d12_instance_RESULT;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_070f4d12_(GO, port_5374d8fd_, RESULT);
input		GO;
input	[15:0]	port_5374d8fd_;
output	[15:0]	RESULT;
wire signed	[15:0]	greaterThan_a_signed;
wire		greaterThan;
wire signed	[15:0]	greaterThan_b_signed;
wire		not_u44_u0;
wire		and_u275_u0;
wire		and_u276_u0;
wire	[15:0]	mux_u20;
wire		and_u277_u0;
wire		and_u278_u0;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_5374d8fd_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign not_u44_u0=~greaterThan;
assign and_u275_u0=GO&greaterThan;
assign and_u276_u0=GO&not_u44_u0;
assign mux_u20=(and_u277_u0)?port_5374d8fd_:16'h0;
assign and_u277_u0=and_u276_u0&GO;
assign and_u278_u0=and_u275_u0&GO;
assign RESULT=mux_u20;
endmodule



module LL1_H_iunzipFilter2D_midNoConsume2(CLK, RESET, GO, port_50b9449e_, port_645796b3_, port_7c5db129_, RESULT, RESULT_u209, RESULT_u210, RESULT_u211, RESULT_u212, RESULT_u213, RESULT_u214, RESULT_u215, RESULT_u216, RESULT_u217, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_50b9449e_;
input		port_645796b3_;
input	[15:0]	port_7c5db129_;
output		RESULT;
output	[15:0]	RESULT_u209;
output		RESULT_u210;
output	[15:0]	RESULT_u211;
output		RESULT_u212;
output	[31:0]	RESULT_u213;
output	[2:0]	RESULT_u214;
output	[15:0]	RESULT_u215;
output	[15:0]	RESULT_u216;
output		RESULT_u217;
output		DONE;
wire		and_u281_u0;
wire		or_u60_u0;
reg		done_cache_u24=1'h0;
reg		done_cache_u25_u0=1'h0;
wire		and_u286_u0;
wire		or_u61_u0;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_0c206b86_instance_RESULT;
wire	[15:0]	add;
wire	[15:0]	simplePinWrite;
wire		simplePinWrite_u56;
wire	[15:0]	simplePinWrite_u57;
reg		reg_492e2661_u0=1'h0;
reg		reg_492e2661_result_delayed_u0=1'h0;
reg	[15:0]	syncEnable_u17=16'h0;
reg		reg_2a40bafa_u0=1'h0;
wire		or_u62_u0;
reg		reg_492e2661_result_delayed_result_delayed_u0=1'h0;
reg		reg_2a40bafa_result_delayed_u0=1'h0;
assign and_u281_u0=done_cache_u24&port_645796b3_;
assign or_u60_u0=and_u281_u0|RESET;
always @(posedge CLK or posedge GO or posedge or_u60_u0)
begin
if (or_u60_u0)
done_cache_u24<=1'h0;
else if (GO)
done_cache_u24<=1'h1;
else done_cache_u24<=done_cache_u24;
end
always @(posedge CLK or posedge reg_2a40bafa_result_delayed_u0 or posedge or_u61_u0)
begin
if (or_u61_u0)
done_cache_u25_u0<=1'h0;
else if (reg_2a40bafa_result_delayed_u0)
done_cache_u25_u0<=1'h1;
else done_cache_u25_u0<=done_cache_u25_u0;
end
assign and_u286_u0=done_cache_u25_u0&port_645796b3_;
assign or_u61_u0=and_u286_u0|RESET;
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_0c206b86_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_0c206b86_instance(.GO(reg_492e2661_u0), 
  .port_4bf8c82c_(syncEnable_u17), .port_4d642370_(port_7c5db129_), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_0c206b86_instance_RESULT));
assign add=port_50b9449e_+16'h1;
assign simplePinWrite=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_0c206b86_instance_RESULT&{16{reg_492e2661_u0}};
assign simplePinWrite_u56=reg_492e2661_u0&{1{reg_492e2661_u0}};
assign simplePinWrite_u57=16'h1&{16{1'h1}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_492e2661_u0<=1'h0;
else reg_492e2661_u0<=reg_2a40bafa_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_492e2661_result_delayed_u0<=1'h0;
else reg_492e2661_result_delayed_u0<=reg_492e2661_u0;
end
always @(posedge CLK)
begin
if (reg_2a40bafa_u0)
syncEnable_u17<=port_7c5db129_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2a40bafa_u0<=1'h0;
else reg_2a40bafa_u0<=GO;
end
assign or_u62_u0=GO|reg_2a40bafa_result_delayed_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_492e2661_result_delayed_result_delayed_u0<=1'h0;
else reg_492e2661_result_delayed_result_delayed_u0<=reg_492e2661_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2a40bafa_result_delayed_u0<=1'h0;
else reg_2a40bafa_result_delayed_u0<=reg_2a40bafa_u0;
end
assign RESULT=GO;
assign RESULT_u209=16'h0;
assign RESULT_u210=GO;
assign RESULT_u211=add;
assign RESULT_u212=or_u62_u0;
assign RESULT_u213=32'h0;
assign RESULT_u214=3'h1;
assign RESULT_u215=simplePinWrite_u57;
assign RESULT_u216=simplePinWrite;
assign RESULT_u217=simplePinWrite_u56;
assign DONE=reg_492e2661_result_delayed_result_delayed_u0;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_0c206b86_(GO, port_4bf8c82c_, port_4d642370_, RESULT);
input		GO;
input	[15:0]	port_4bf8c82c_;
input	[15:0]	port_4d642370_;
output	[15:0]	RESULT;
wire	[15:0]	subtract;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_5f781e45_instance_RESULT;
assign subtract=port_4bf8c82c_-port_4d642370_;
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_5f781e45_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_5f781e45_instance(.GO(GO), 
  .port_399b2cce_({subtract[15], subtract[15:1]}), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_5f781e45_instance_RESULT));
assign RESULT=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_5f781e45_instance_RESULT;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_5f781e45_(GO, port_399b2cce_, RESULT);
input		GO;
input	[15:0]	port_399b2cce_;
output	[15:0]	RESULT;
wire signed	[15:0]	greaterThan_b_signed;
wire		greaterThan;
wire signed	[15:0]	greaterThan_a_signed;
wire		and_u290_u0;
wire		and_u291_u0;
wire		not_u45_u0;
wire		and_u292_u0;
wire		and_u293_u0;
wire	[15:0]	mux_u21;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_399b2cce_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign and_u290_u0=GO&greaterThan;
assign and_u291_u0=GO&not_u45_u0;
assign not_u45_u0=~greaterThan;
assign and_u292_u0=and_u290_u0&GO;
assign and_u293_u0=and_u291_u0&GO;
assign mux_u21=(and_u293_u0)?port_399b2cce_:16'h0;
assign RESULT=mux_u21;
endmodule



module LL1_H_iunzipFilter2D_simplememoryreferee_6b7a23db_(bus_5baae8ff_, bus_7653fefb_, bus_341c19c0_, bus_31af2b27_, bus_3c374e45_, bus_6913617c_, bus_2cde6fec_, bus_3374a16b_, bus_19f443bd_, bus_1553ab35_, bus_663891ac_, bus_15e55fff_, bus_0d5861d7_, bus_53cfd8c7_, bus_597c15fe_, bus_5900c238_, bus_524805ba_, bus_3a1a33d5_, bus_3c586cf4_, bus_3c30ecac_, bus_572c858a_, bus_75f74205_, bus_38f192ff_, bus_675a6465_, bus_4185e507_, bus_38250251_, bus_03b2b05f_, bus_7654652b_, bus_51b62008_, bus_5930e896_, bus_182c3189_, bus_472d9480_, bus_1ec5415f_, bus_1291fb88_, bus_0a2e3320_, bus_72eea4ff_, bus_77976b59_, bus_3af85b4e_, bus_499884d1_, bus_1b25f6ba_, bus_74cb0e55_, bus_756e636f_, bus_06803267_, bus_02376507_, bus_3be386e2_, bus_013e7d74_, bus_37e5e149_, bus_0512548f_, bus_398aca9c_, bus_007ee040_, bus_1d49e0c0_, bus_1c6c6256_, bus_08b6bf94_, bus_06d6df27_, bus_74b6e615_, bus_63d1ee63_, bus_2a8034ec_, bus_597f939d_, bus_309722e6_, bus_783c1160_, bus_3295fff5_, bus_66b8fa73_, bus_27bf1f93_, bus_56c466b1_, bus_3ab47106_, bus_562d02e1_, bus_194c7c11_, bus_68a5f92c_, bus_3fe7f593_, bus_3c0153f0_, bus_22677e1d_, bus_0fc79387_, bus_55cc71ee_, bus_084108ff_, bus_60937d22_, bus_39138d0a_, bus_38f0c907_, bus_1be8460e_, bus_546e4ea1_, bus_68c80959_, bus_723f4da1_, bus_118dcb12_, bus_34e6dfec_, bus_47803ec7_, bus_5eb5ed16_, bus_1807f3cd_, bus_1446f926_, bus_7b461753_, bus_1df60b90_, bus_4ad1a98a_, bus_7b6d2db0_, bus_295fc32e_, bus_42424c02_, bus_05553665_, bus_75b6e6aa_, bus_782a49ae_, bus_167da5bd_, bus_7e378a50_, bus_03a2926d_, bus_299c5c34_, bus_12066278_, bus_31710b5f_, bus_27d78a2b_, bus_78fb14d7_, bus_52935bd9_, bus_5122026c_, bus_35bb43c2_, bus_1f5c5926_, bus_7cd6911c_, bus_57083dd4_, bus_2f7aa6e4_, bus_0ad99597_, bus_5a5f2961_, bus_2781fc25_, bus_02c8854d_, bus_3b77c854_, bus_6308ab98_, bus_78addd53_, bus_2c656446_, bus_15fa8b31_, bus_29c7540a_, bus_24ac86a8_, bus_623e353f_, bus_0fd98caa_, bus_4b3e6981_, bus_75734968_, bus_5727ff78_, bus_018f435a_, bus_13a61289_, bus_6341aa95_, bus_5a1ddee7_, bus_47b6d4cf_);
input		bus_5baae8ff_;
input		bus_7653fefb_;
input		bus_341c19c0_;
input	[15:0]	bus_31af2b27_;
input		bus_3c374e45_;
input		bus_6913617c_;
input	[15:0]	bus_2cde6fec_;
input	[31:0]	bus_3374a16b_;
input	[2:0]	bus_19f443bd_;
input		bus_1553ab35_;
input		bus_663891ac_;
input	[15:0]	bus_15e55fff_;
input	[31:0]	bus_0d5861d7_;
input	[2:0]	bus_53cfd8c7_;
input		bus_597c15fe_;
input		bus_5900c238_;
input	[15:0]	bus_524805ba_;
input	[31:0]	bus_3a1a33d5_;
input	[2:0]	bus_3c586cf4_;
input		bus_3c30ecac_;
input		bus_572c858a_;
input	[15:0]	bus_75f74205_;
input	[31:0]	bus_38f192ff_;
input	[2:0]	bus_675a6465_;
input		bus_4185e507_;
input		bus_38250251_;
input	[15:0]	bus_03b2b05f_;
input	[31:0]	bus_7654652b_;
input	[2:0]	bus_51b62008_;
input		bus_5930e896_;
input	[31:0]	bus_182c3189_;
input	[2:0]	bus_472d9480_;
input		bus_1ec5415f_;
input	[31:0]	bus_1291fb88_;
input	[2:0]	bus_0a2e3320_;
input		bus_72eea4ff_;
input		bus_77976b59_;
input	[15:0]	bus_3af85b4e_;
input	[31:0]	bus_499884d1_;
input	[2:0]	bus_1b25f6ba_;
input		bus_74cb0e55_;
input		bus_756e636f_;
input	[15:0]	bus_06803267_;
input	[31:0]	bus_02376507_;
input	[2:0]	bus_3be386e2_;
input		bus_013e7d74_;
input	[31:0]	bus_37e5e149_;
input	[2:0]	bus_0512548f_;
input		bus_398aca9c_;
input	[31:0]	bus_007ee040_;
input	[2:0]	bus_1d49e0c0_;
input		bus_1c6c6256_;
input		bus_08b6bf94_;
input	[15:0]	bus_06d6df27_;
input	[31:0]	bus_74b6e615_;
input	[2:0]	bus_63d1ee63_;
input		bus_2a8034ec_;
input		bus_597f939d_;
input	[15:0]	bus_309722e6_;
input	[31:0]	bus_783c1160_;
input	[2:0]	bus_3295fff5_;
input		bus_66b8fa73_;
input	[31:0]	bus_27bf1f93_;
input	[2:0]	bus_56c466b1_;
input		bus_3ab47106_;
input	[31:0]	bus_562d02e1_;
input	[2:0]	bus_194c7c11_;
input		bus_68a5f92c_;
input	[31:0]	bus_3fe7f593_;
input	[2:0]	bus_3c0153f0_;
input		bus_22677e1d_;
input	[31:0]	bus_0fc79387_;
input	[2:0]	bus_55cc71ee_;
input		bus_084108ff_;
input	[31:0]	bus_60937d22_;
input	[2:0]	bus_39138d0a_;
input		bus_38f0c907_;
input	[31:0]	bus_1be8460e_;
input	[2:0]	bus_546e4ea1_;
input		bus_68c80959_;
input	[31:0]	bus_723f4da1_;
input	[2:0]	bus_118dcb12_;
input		bus_34e6dfec_;
input	[31:0]	bus_47803ec7_;
input	[2:0]	bus_5eb5ed16_;
output	[15:0]	bus_1807f3cd_;
output	[31:0]	bus_1446f926_;
output		bus_7b461753_;
output		bus_1df60b90_;
output	[2:0]	bus_4ad1a98a_;
output	[15:0]	bus_7b6d2db0_;
output		bus_295fc32e_;
output	[15:0]	bus_42424c02_;
output		bus_05553665_;
output	[15:0]	bus_75b6e6aa_;
output		bus_782a49ae_;
output	[15:0]	bus_167da5bd_;
output		bus_7e378a50_;
output	[15:0]	bus_03a2926d_;
output		bus_299c5c34_;
output	[15:0]	bus_12066278_;
output		bus_31710b5f_;
output	[15:0]	bus_27d78a2b_;
output		bus_78fb14d7_;
output	[15:0]	bus_52935bd9_;
output		bus_5122026c_;
output	[15:0]	bus_35bb43c2_;
output		bus_1f5c5926_;
output	[15:0]	bus_7cd6911c_;
output		bus_57083dd4_;
output	[15:0]	bus_2f7aa6e4_;
output		bus_0ad99597_;
output	[15:0]	bus_5a5f2961_;
output		bus_2781fc25_;
output	[15:0]	bus_02c8854d_;
output		bus_3b77c854_;
output	[15:0]	bus_6308ab98_;
output		bus_78addd53_;
output	[15:0]	bus_2c656446_;
output		bus_15fa8b31_;
output	[15:0]	bus_29c7540a_;
output		bus_24ac86a8_;
output	[15:0]	bus_623e353f_;
output		bus_0fd98caa_;
output	[15:0]	bus_4b3e6981_;
output		bus_75734968_;
output	[15:0]	bus_5727ff78_;
output		bus_018f435a_;
output	[15:0]	bus_13a61289_;
output		bus_6341aa95_;
output	[15:0]	bus_5a1ddee7_;
output		bus_47b6d4cf_;
wire		or_173d943c_u0;
wire		not_5ea54ea7_u0;
wire		or_1129842a_u0;
wire		not_6ad8d1dd_u0;
wire		and_787f997a_u0;
wire		not_4e7f7c71_u0;
reg		done_qual_u0=1'h0;
wire		not_26eb2efb_u0;
reg		done_qual_u1_u0=1'h0;
wire		and_50ece2f9_u0;
reg		done_qual_u2_u0=1'h0;
wire		or_1675ff6c_u0;
wire		not_4746555d_u0;
reg		done_qual_u3_u0=1'h0;
wire		not_0ea8a9b6_u0;
wire		not_17a0b380_u0;
reg		done_qual_u4_u0=1'h0;
reg		done_qual_u5_u0=1'h0;
wire		or_3c053826_u0;
wire		and_1cf374d4_u0;
wire		or_1f537b7b_u0;
wire		and_730e8f24_u0;
reg		done_qual_u6_u0=1'h0;
wire		or_4d04e829_u0;
wire		or_733bc914_u0;
wire		or_6b0d213c_u0;
wire		and_150a423f_u0;
wire		not_12465171_u0;
wire		or_663a9602_u0;
wire		not_2c5be261_u0;
wire		or_41aa7f90_u0;
wire		or_6b55ce68_u0;
wire		not_2e950ad6_u0;
wire		not_2d18c45e_u0;
wire		or_3e8674c1_u0;
reg		done_qual_u7_u0=1'h0;
reg		done_qual_u8_u0=1'h0;
wire		not_2abc77ed_u0;
wire		not_3cf708a6_u0;
reg		done_qual_u9_u0=1'h0;
wire		not_349670c0_u0;
wire		or_5ac66791_u0;
wire		and_5f9d39c1_u0;
wire		and_36c210a0_u0;
wire		and_35511b36_u0;
wire		or_15a163c9_u0;
wire		and_3de7018d_u0;
wire		and_702a8b40_u0;
reg		done_qual_u10_u0=1'h0;
reg		done_qual_u11_u0=1'h0;
wire		or_2b55e325_u0;
reg		done_qual_u12_u0=1'h0;
wire		and_209011e4_u0;
wire		or_12432836_u0;
wire		or_3e44203e_u0;
wire		or_5f6d6716_u0;
wire		or_5e493e35_u0;
wire		or_4add4d5f_u0;
wire		or_1f7711f0_u0;
wire		and_3fccd641_u0;
wire		or_1633f2a1_u0;
wire		or_08eb4378_u0;
wire		not_70d80b4d_u0;
reg		done_qual_u13_u0=1'h0;
wire		and_175b1ec3_u0;
wire		or_0b06549a_u0;
reg		done_qual_u14_u0=1'h0;
reg		done_qual_u15_u0=1'h0;
wire		or_05e1be52_u0;
wire		not_60a2b111_u0;
wire		and_0508babc_u0;
wire		and_75df8e69_u0;
reg		done_qual_u16_u0=1'h0;
wire	[31:0]	mux_1be6495d_u0;
reg		done_qual_u17_u0=1'h0;
reg		done_qual_u18_u0=1'h0;
wire		not_73ce8707_u0;
wire		and_0d6698ac_u0;
wire		and_7a892d46_u0;
wire		or_69a9fb7a_u0;
wire		not_7f8b7458_u0;
wire		or_7cf5ad22_u0;
wire		or_1f3cbcdd_u0;
wire		or_4f4e3ba6_u0;
wire		or_10e5e40d_u0;
reg		done_qual_u19_u0=1'h0;
wire		or_562e18df_u0;
wire		and_154ea8b9_u0;
reg		done_qual_u20_u0=1'h0;
wire		and_0319b9ee_u0;
wire		not_5bcead36_u0;
wire		and_68495db0_u0;
wire		not_6426c4dd_u0;
wire		and_76f7b10c_u0;
wire		not_6c9ef860_u0;
wire	[15:0]	mux_038b2974_u0;
wire		or_66865279_u0;
assign or_173d943c_u0=bus_3c30ecac_|bus_572c858a_;
assign not_5ea54ea7_u0=~bus_341c19c0_;
assign or_1129842a_u0=or_3e8674c1_u0|done_qual_u15_u0;
assign not_6ad8d1dd_u0=~bus_341c19c0_;
assign and_787f997a_u0=or_1675ff6c_u0&bus_341c19c0_;
assign not_4e7f7c71_u0=~bus_341c19c0_;
always @(posedge bus_5baae8ff_)
begin
if (bus_7653fefb_)
done_qual_u0<=1'h0;
else done_qual_u0<=bus_084108ff_;
end
assign not_26eb2efb_u0=~bus_341c19c0_;
always @(posedge bus_5baae8ff_)
begin
if (bus_7653fefb_)
done_qual_u1_u0<=1'h0;
else done_qual_u1_u0<=bus_3ab47106_;
end
assign and_50ece2f9_u0=or_4f4e3ba6_u0&bus_341c19c0_;
always @(posedge bus_5baae8ff_)
begin
if (bus_7653fefb_)
done_qual_u2_u0<=1'h0;
else done_qual_u2_u0<=or_3e44203e_u0;
end
assign or_1675ff6c_u0=or_733bc914_u0|done_qual_u7_u0;
assign not_4746555d_u0=~bus_341c19c0_;
always @(posedge bus_5baae8ff_)
begin
if (bus_7653fefb_)
done_qual_u3_u0<=1'h0;
else done_qual_u3_u0<=or_173d943c_u0;
end
assign not_0ea8a9b6_u0=~bus_341c19c0_;
assign not_17a0b380_u0=~bus_341c19c0_;
always @(posedge bus_5baae8ff_)
begin
if (bus_7653fefb_)
done_qual_u4_u0<=1'h0;
else done_qual_u4_u0<=bus_013e7d74_;
end
always @(posedge bus_5baae8ff_)
begin
if (bus_7653fefb_)
done_qual_u5_u0<=1'h0;
else done_qual_u5_u0<=or_1f7711f0_u0;
end
assign or_3c053826_u0=bus_34e6dfec_|done_qual_u9_u0;
assign and_1cf374d4_u0=or_15a163c9_u0&bus_341c19c0_;
assign or_1f537b7b_u0=or_41aa7f90_u0|done_qual_u19_u0;
assign and_730e8f24_u0=or_4d04e829_u0&bus_341c19c0_;
always @(posedge bus_5baae8ff_)
begin
if (bus_7653fefb_)
done_qual_u6_u0<=1'h0;
else done_qual_u6_u0<=bus_66b8fa73_;
end
assign or_4d04e829_u0=bus_3ab47106_|done_qual_u1_u0;
assign or_733bc914_u0=bus_72eea4ff_|bus_77976b59_;
assign or_6b0d213c_u0=bus_2a8034ec_|bus_597f939d_;
assign and_150a423f_u0=or_663a9602_u0&bus_341c19c0_;
assign not_12465171_u0=~bus_341c19c0_;
assign or_663a9602_u0=or_6b0d213c_u0|done_qual_u10_u0;
assign not_2c5be261_u0=~bus_341c19c0_;
assign or_41aa7f90_u0=bus_4185e507_|bus_38250251_;
assign or_6b55ce68_u0=bus_6913617c_|bus_663891ac_|bus_5900c238_|bus_572c858a_|bus_38250251_|bus_77976b59_|bus_756e636f_|bus_08b6bf94_|bus_597f939d_;
assign not_2e950ad6_u0=~bus_341c19c0_;
assign not_2d18c45e_u0=~bus_341c19c0_;
assign or_3e8674c1_u0=bus_597c15fe_|bus_5900c238_;
always @(posedge bus_5baae8ff_)
begin
if (bus_7653fefb_)
done_qual_u7_u0<=1'h0;
else done_qual_u7_u0<=or_733bc914_u0;
end
assign bus_1807f3cd_=mux_038b2974_u0;
assign bus_1446f926_=mux_1be6495d_u0;
assign bus_7b461753_=or_6b55ce68_u0;
assign bus_1df60b90_=or_1633f2a1_u0;
assign bus_4ad1a98a_=3'h1;
assign bus_7b6d2db0_=bus_31af2b27_;
assign bus_295fc32e_=and_1cf374d4_u0;
assign bus_42424c02_=bus_31af2b27_;
assign bus_05553665_=and_209011e4_u0;
assign bus_75b6e6aa_=bus_31af2b27_;
assign bus_782a49ae_=and_7a892d46_u0;
assign bus_167da5bd_=bus_31af2b27_;
assign bus_7e378a50_=and_175b1ec3_u0;
assign bus_03a2926d_=bus_31af2b27_;
assign bus_299c5c34_=and_0d6698ac_u0;
assign bus_12066278_=bus_31af2b27_;
assign bus_31710b5f_=and_35511b36_u0;
assign bus_27d78a2b_=bus_31af2b27_;
assign bus_78fb14d7_=and_36c210a0_u0;
assign bus_52935bd9_=bus_31af2b27_;
assign bus_5122026c_=and_787f997a_u0;
assign bus_35bb43c2_=bus_31af2b27_;
assign bus_1f5c5926_=and_76f7b10c_u0;
assign bus_7cd6911c_=bus_31af2b27_;
assign bus_57083dd4_=and_50ece2f9_u0;
assign bus_2f7aa6e4_=bus_31af2b27_;
assign bus_0ad99597_=and_68495db0_u0;
assign bus_5a5f2961_=bus_31af2b27_;
assign bus_2781fc25_=and_5f9d39c1_u0;
assign bus_02c8854d_=bus_31af2b27_;
assign bus_3b77c854_=and_150a423f_u0;
assign bus_6308ab98_=bus_31af2b27_;
assign bus_78addd53_=and_154ea8b9_u0;
assign bus_2c656446_=bus_31af2b27_;
assign bus_15fa8b31_=and_730e8f24_u0;
assign bus_29c7540a_=bus_31af2b27_;
assign bus_24ac86a8_=and_75df8e69_u0;
assign bus_623e353f_=bus_31af2b27_;
assign bus_0fd98caa_=and_3de7018d_u0;
assign bus_4b3e6981_=bus_31af2b27_;
assign bus_75734968_=and_0508babc_u0;
assign bus_5727ff78_=bus_31af2b27_;
assign bus_018f435a_=and_0319b9ee_u0;
assign bus_13a61289_=bus_31af2b27_;
assign bus_6341aa95_=and_702a8b40_u0;
assign bus_5a1ddee7_=bus_31af2b27_;
assign bus_47b6d4cf_=and_3fccd641_u0;
always @(posedge bus_5baae8ff_)
begin
if (bus_7653fefb_)
done_qual_u8_u0<=1'h0;
else done_qual_u8_u0<=bus_5930e896_;
end
assign not_2abc77ed_u0=~bus_341c19c0_;
assign not_3cf708a6_u0=~bus_341c19c0_;
always @(posedge bus_5baae8ff_)
begin
if (bus_7653fefb_)
done_qual_u9_u0<=1'h0;
else done_qual_u9_u0<=bus_34e6dfec_;
end
assign not_349670c0_u0=~bus_341c19c0_;
assign or_5ac66791_u0=bus_22677e1d_|done_qual_u17_u0;
assign and_5f9d39c1_u0=or_1f3cbcdd_u0&bus_341c19c0_;
assign and_36c210a0_u0=or_12432836_u0&bus_341c19c0_;
assign and_35511b36_u0=or_2b55e325_u0&bus_341c19c0_;
assign or_15a163c9_u0=or_69a9fb7a_u0|done_qual_u16_u0;
assign and_3de7018d_u0=or_5ac66791_u0&bus_341c19c0_;
assign and_702a8b40_u0=or_10e5e40d_u0&bus_341c19c0_;
always @(posedge bus_5baae8ff_)
begin
if (bus_7653fefb_)
done_qual_u10_u0<=1'h0;
else done_qual_u10_u0<=or_6b0d213c_u0;
end
always @(posedge bus_5baae8ff_)
begin
if (bus_7653fefb_)
done_qual_u11_u0<=1'h0;
else done_qual_u11_u0<=bus_68a5f92c_;
end
assign or_2b55e325_u0=bus_5930e896_|done_qual_u8_u0;
always @(posedge bus_5baae8ff_)
begin
if (bus_7653fefb_)
done_qual_u12_u0<=1'h0;
else done_qual_u12_u0<=bus_1ec5415f_;
end
assign and_209011e4_u0=or_05e1be52_u0&bus_341c19c0_;
assign or_12432836_u0=bus_1ec5415f_|done_qual_u12_u0;
assign or_3e44203e_u0=bus_1c6c6256_|bus_08b6bf94_;
assign or_5f6d6716_u0=bus_38f0c907_|done_qual_u20_u0;
assign or_5e493e35_u0=bus_66b8fa73_|done_qual_u6_u0;
assign or_4add4d5f_u0=or_173d943c_u0|done_qual_u3_u0;
assign or_1f7711f0_u0=bus_74cb0e55_|bus_756e636f_;
assign and_3fccd641_u0=or_3c053826_u0&bus_341c19c0_;
assign or_1633f2a1_u0=or_69a9fb7a_u0|or_562e18df_u0|or_3e8674c1_u0|or_173d943c_u0|or_41aa7f90_u0|bus_5930e896_|bus_1ec5415f_|or_733bc914_u0|or_1f7711f0_u0|bus_013e7d74_|bus_398aca9c_|or_3e44203e_u0|or_6b0d213c_u0|bus_66b8fa73_|bus_3ab47106_|bus_68a5f92c_|bus_22677e1d_|bus_084108ff_|bus_38f0c907_|bus_68c80959_|bus_34e6dfec_;
assign or_08eb4378_u0=bus_084108ff_|done_qual_u0;
assign not_70d80b4d_u0=~bus_341c19c0_;
always @(posedge bus_5baae8ff_)
begin
if (bus_7653fefb_)
done_qual_u13_u0<=1'h0;
else done_qual_u13_u0<=or_562e18df_u0;
end
assign and_175b1ec3_u0=or_4add4d5f_u0&bus_341c19c0_;
assign or_0b06549a_u0=or_1f7711f0_u0|done_qual_u5_u0;
always @(posedge bus_5baae8ff_)
begin
if (bus_7653fefb_)
done_qual_u14_u0<=1'h0;
else done_qual_u14_u0<=bus_68c80959_;
end
always @(posedge bus_5baae8ff_)
begin
if (bus_7653fefb_)
done_qual_u15_u0<=1'h0;
else done_qual_u15_u0<=or_3e8674c1_u0;
end
assign or_05e1be52_u0=or_562e18df_u0|done_qual_u13_u0;
assign not_60a2b111_u0=~bus_341c19c0_;
assign and_0508babc_u0=or_08eb4378_u0&bus_341c19c0_;
assign and_75df8e69_u0=or_7cf5ad22_u0&bus_341c19c0_;
always @(posedge bus_5baae8ff_)
begin
if (bus_7653fefb_)
done_qual_u16_u0<=1'h0;
else done_qual_u16_u0<=or_69a9fb7a_u0;
end
assign mux_1be6495d_u0=({32{or_69a9fb7a_u0}}&bus_3374a16b_)|({32{or_562e18df_u0}}&32'h0)|({32{or_3e8674c1_u0}}&32'h0)|({32{or_173d943c_u0}}&32'h0)|({32{or_41aa7f90_u0}}&32'h0)|({32{bus_5930e896_}}&32'h0)|({32{bus_1ec5415f_}}&32'h0)|({32{or_733bc914_u0}}&32'h0)|({32{or_1f7711f0_u0}}&32'h0)|({32{bus_013e7d74_}}&32'h0)|({32{bus_398aca9c_}}&32'h0)|({32{or_3e44203e_u0}}&32'h0)|({32{or_6b0d213c_u0}}&32'h0)|({32{bus_66b8fa73_}}&32'h0)|({32{bus_3ab47106_}}&32'h0)|({32{bus_68a5f92c_}}&32'h0)|({32{bus_22677e1d_}}&32'h0)|({32{bus_084108ff_}}&32'h0)|({32{bus_38f0c907_}}&32'h0)|({32{bus_68c80959_}}&32'h0)|({32{bus_34e6dfec_}}&32'h0);
always @(posedge bus_5baae8ff_)
begin
if (bus_7653fefb_)
done_qual_u17_u0<=1'h0;
else done_qual_u17_u0<=bus_22677e1d_;
end
always @(posedge bus_5baae8ff_)
begin
if (bus_7653fefb_)
done_qual_u18_u0<=1'h0;
else done_qual_u18_u0<=bus_398aca9c_;
end
assign not_73ce8707_u0=~bus_341c19c0_;
assign and_0d6698ac_u0=or_1f537b7b_u0&bus_341c19c0_;
assign and_7a892d46_u0=or_1129842a_u0&bus_341c19c0_;
assign or_69a9fb7a_u0=bus_3c374e45_|bus_6913617c_;
assign not_7f8b7458_u0=~bus_341c19c0_;
assign or_7cf5ad22_u0=bus_68a5f92c_|done_qual_u11_u0;
assign or_1f3cbcdd_u0=or_3e44203e_u0|done_qual_u2_u0;
assign or_4f4e3ba6_u0=bus_013e7d74_|done_qual_u4_u0;
assign or_10e5e40d_u0=bus_68c80959_|done_qual_u14_u0;
always @(posedge bus_5baae8ff_)
begin
if (bus_7653fefb_)
done_qual_u19_u0<=1'h0;
else done_qual_u19_u0<=or_41aa7f90_u0;
end
assign or_562e18df_u0=bus_1553ab35_|bus_663891ac_;
assign and_154ea8b9_u0=or_5e493e35_u0&bus_341c19c0_;
always @(posedge bus_5baae8ff_)
begin
if (bus_7653fefb_)
done_qual_u20_u0<=1'h0;
else done_qual_u20_u0<=bus_38f0c907_;
end
assign and_0319b9ee_u0=or_5f6d6716_u0&bus_341c19c0_;
assign not_5bcead36_u0=~bus_341c19c0_;
assign and_68495db0_u0=or_66865279_u0&bus_341c19c0_;
assign not_6426c4dd_u0=~bus_341c19c0_;
assign and_76f7b10c_u0=or_0b06549a_u0&bus_341c19c0_;
assign not_6c9ef860_u0=~bus_341c19c0_;
assign mux_038b2974_u0=({16{bus_6913617c_}}&bus_2cde6fec_)|({16{bus_663891ac_}}&bus_15e55fff_)|({16{bus_5900c238_}}&bus_524805ba_)|({16{bus_572c858a_}}&bus_75f74205_)|({16{bus_38250251_}}&bus_03b2b05f_)|({16{bus_77976b59_}}&bus_3af85b4e_)|({16{bus_756e636f_}}&bus_06803267_)|({16{bus_08b6bf94_}}&bus_06d6df27_)|({16{bus_597f939d_}}&bus_309722e6_);
assign or_66865279_u0=bus_398aca9c_|done_qual_u18_u0;
endmodule



module LL1_H_iunzipFilter2D_topRow(CLK, RESET, GO, port_72b95caa_, port_43ed3c0e_, port_3b2ce771_, port_758e77d7_, port_0b4ae4bc_, port_59b37350_, port_054c182e_, RESULT, RESULT_u218, RESULT_u219, RESULT_u220, RESULT_u221, RESULT_u222, RESULT_u223, RESULT_u224, RESULT_u225, RESULT_u226, RESULT_u227, RESULT_u228, RESULT_u229, RESULT_u230, RESULT_u231, RESULT_u232, RESULT_u233, RESULT_u234, RESULT_u235, DONE);
input		CLK;
input		RESET;
input		GO;
input	[31:0]	port_72b95caa_;
input	[15:0]	port_43ed3c0e_;
input	[15:0]	port_3b2ce771_;
input		port_758e77d7_;
input	[15:0]	port_0b4ae4bc_;
input		port_59b37350_;
input	[15:0]	port_054c182e_;
output		RESULT;
output	[31:0]	RESULT_u218;
output		RESULT_u219;
output	[15:0]	RESULT_u220;
output		RESULT_u221;
output	[15:0]	RESULT_u222;
output		RESULT_u223;
output	[15:0]	RESULT_u224;
output		RESULT_u225;
output	[31:0]	RESULT_u226;
output	[2:0]	RESULT_u227;
output		RESULT_u228;
output	[31:0]	RESULT_u229;
output	[15:0]	RESULT_u230;
output	[2:0]	RESULT_u231;
output		RESULT_u232;
output	[15:0]	RESULT_u233;
output		RESULT_u234;
output	[15:0]	RESULT_u235;
output		DONE;
wire		simplePinWrite;
wire		and_u296_u0;
wire		or_u63_u0;
reg		done_cache_u26=1'h0;
wire		or_u64_u0;
reg		done_cache_u27_u0=1'h0;
wire		and_u300_u0;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_2459cdf0_instance_RESULT;
reg		reg_59bcaa5a_u0=1'h0;
wire		and_u309_u0;
wire		or_u65_u0;
wire	[31:0]	add;
wire	[15:0]	add_u4;
wire	[15:0]	add_u5;
wire		simplePinWrite_u58;
wire	[15:0]	simplePinWrite_u59;
wire	[15:0]	simplePinWrite_u60;
reg		reg_575a9c62_u0=1'h0;
wire		or_u66_u0;
reg		reg_27cfe5ac_u0=1'h0;
reg		reg_6546ce30_u0=1'h0;
reg		reg_575a9c62_result_delayed_u0=1'h0;
reg		reg_28c7b954_u0=1'h0;
reg	[15:0]	syncEnable_u18=16'h0;
reg		reg_6546ce30_result_delayed_u0=1'h0;
reg	[15:0]	syncEnable_u19_u0=16'h0;
assign simplePinWrite=GO&{1{GO}};
assign and_u296_u0=done_cache_u26&port_59b37350_;
assign or_u63_u0=and_u296_u0|RESET;
always @(posedge CLK or posedge GO or posedge or_u63_u0)
begin
if (or_u63_u0)
done_cache_u26<=1'h0;
else if (GO)
done_cache_u26<=1'h1;
else done_cache_u26<=done_cache_u26;
end
assign or_u64_u0=and_u300_u0|RESET;
always @(posedge CLK or posedge reg_6546ce30_result_delayed_u0 or posedge or_u64_u0)
begin
if (or_u64_u0)
done_cache_u27_u0<=1'h0;
else if (reg_6546ce30_result_delayed_u0)
done_cache_u27_u0<=1'h1;
else done_cache_u27_u0<=done_cache_u27_u0;
end
assign and_u300_u0=done_cache_u27_u0&port_59b37350_;
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_2459cdf0_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_2459cdf0_instance(.GO(reg_28c7b954_u0), 
  .port_6f393820_(port_0b4ae4bc_), .port_40d4a25f_(syncEnable_u18), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_2459cdf0_instance_RESULT));
always @(posedge CLK or posedge reg_575a9c62_result_delayed_u0 or posedge or_u65_u0)
begin
if (or_u65_u0)
reg_59bcaa5a_u0<=1'h0;
else if (reg_575a9c62_result_delayed_u0)
reg_59bcaa5a_u0<=1'h1;
else reg_59bcaa5a_u0<=reg_59bcaa5a_u0;
end
assign and_u309_u0=reg_59bcaa5a_u0&port_59b37350_;
assign or_u65_u0=and_u309_u0|RESET;
assign add=port_72b95caa_+32'h1;
assign add_u4=port_43ed3c0e_+16'h1;
assign add_u5=port_3b2ce771_+16'h1;
assign simplePinWrite_u58=reg_28c7b954_u0&{1{reg_28c7b954_u0}};
assign simplePinWrite_u59=16'h1&{16{1'h1}};
assign simplePinWrite_u60=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_2459cdf0_instance_RESULT&{16{reg_28c7b954_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_575a9c62_u0<=1'h0;
else reg_575a9c62_u0<=reg_28c7b954_u0;
end
assign or_u66_u0=GO|reg_6546ce30_result_delayed_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_27cfe5ac_u0<=1'h0;
else reg_27cfe5ac_u0<=reg_575a9c62_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6546ce30_u0<=1'h0;
else reg_6546ce30_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_575a9c62_result_delayed_u0<=1'h0;
else reg_575a9c62_result_delayed_u0<=reg_575a9c62_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_28c7b954_u0<=1'h0;
else reg_28c7b954_u0<=reg_6546ce30_result_delayed_u0;
end
always @(posedge CLK)
begin
if (reg_6546ce30_u0)
syncEnable_u18<=port_0b4ae4bc_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6546ce30_result_delayed_u0<=1'h0;
else reg_6546ce30_result_delayed_u0<=reg_6546ce30_u0;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u19_u0<=port_054c182e_;
end
assign RESULT=GO;
assign RESULT_u218=add;
assign RESULT_u219=GO;
assign RESULT_u220=16'h0;
assign RESULT_u221=GO;
assign RESULT_u222=add_u4;
assign RESULT_u223=GO;
assign RESULT_u224=add_u5;
assign RESULT_u225=or_u66_u0;
assign RESULT_u226=32'h0;
assign RESULT_u227=3'h1;
assign RESULT_u228=reg_575a9c62_result_delayed_u0;
assign RESULT_u229=32'h0;
assign RESULT_u230=syncEnable_u19_u0;
assign RESULT_u231=3'h1;
assign RESULT_u232=simplePinWrite;
assign RESULT_u233=simplePinWrite_u59;
assign RESULT_u234=simplePinWrite_u58;
assign RESULT_u235=simplePinWrite_u60;
assign DONE=reg_27cfe5ac_u0;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_2459cdf0_(GO, port_6f393820_, port_40d4a25f_, RESULT);
input		GO;
input	[15:0]	port_6f393820_;
input	[15:0]	port_40d4a25f_;
output	[15:0]	RESULT;
wire	[16:0]	add;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_11e9a72f_instance_RESULT;
assign add={port_40d4a25f_[15], port_40d4a25f_}+{port_6f393820_[15], port_6f393820_};
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_11e9a72f_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_11e9a72f_instance(.GO(GO), 
  .port_0ae41dc7_({add[16], add[16:2]}), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_11e9a72f_instance_RESULT));
assign RESULT=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_11e9a72f_instance_RESULT;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_11e9a72f_(GO, port_0ae41dc7_, RESULT);
input		GO;
input	[15:0]	port_0ae41dc7_;
output	[15:0]	RESULT;
wire signed	[15:0]	greaterThan_b_signed;
wire		greaterThan;
wire signed	[15:0]	greaterThan_a_signed;
wire		not_u46_u0;
wire		and_u304_u0;
wire		and_u305_u0;
wire		and_u306_u0;
wire	[15:0]	mux_u22;
wire		and_u307_u0;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_0ae41dc7_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign not_u46_u0=~greaterThan;
assign and_u304_u0=GO&not_u46_u0;
assign and_u305_u0=GO&greaterThan;
assign and_u306_u0=and_u304_u0&GO;
assign mux_u22=(and_u307_u0)?16'h0:port_0ae41dc7_;
assign and_u307_u0=and_u305_u0&GO;
assign RESULT=mux_u22;
endmodule



module LL1_H_iunzipFilter2D_endianswapper_077bd2d3_(endianswapper_077bd2d3_in, endianswapper_077bd2d3_out);
input	[15:0]	endianswapper_077bd2d3_in;
output	[15:0]	endianswapper_077bd2d3_out;
assign endianswapper_077bd2d3_out=16'h0;
endmodule



module LL1_H_iunzipFilter2D_endianswapper_6f898fe2_(endianswapper_6f898fe2_in, endianswapper_6f898fe2_out);
input	[15:0]	endianswapper_6f898fe2_in;
output	[15:0]	endianswapper_6f898fe2_out;
assign endianswapper_6f898fe2_out=16'h0;
endmodule



module LL1_H_iunzipFilter2D_stateVar_idx(bus_0cf2d3f5_, bus_068d6c06_, bus_674bf37e_, bus_10bc57e4_, bus_4a2d20e1_, bus_22b29207_, bus_5c4dede9_, bus_253147b9_, bus_4ebaa98e_, bus_5ceaaebb_, bus_63833c02_, bus_50790775_, bus_2264995f_, bus_1cdbfe01_, bus_2c539ca8_, bus_632c90cd_, bus_2397b779_, bus_26b5b1f6_, bus_2570bc16_, bus_48005bbe_, bus_441deb71_, bus_46b2645c_, bus_62a23944_, bus_1378e939_, bus_513697cc_, bus_2cee4380_, bus_0475cc13_, bus_78940204_, bus_766fd037_, bus_4d505dca_, bus_1de90dae_, bus_20ace7e3_, bus_1c515fcc_, bus_5e13118c_, bus_041f2681_, bus_6056c028_, bus_3aa04241_, bus_3321cb07_, bus_7e50ec6c_, bus_26d18263_, bus_2a7d4abb_);
input		bus_0cf2d3f5_;
input		bus_068d6c06_;
input		bus_674bf37e_;
input	[15:0]	bus_10bc57e4_;
input		bus_4a2d20e1_;
input	[15:0]	bus_22b29207_;
input		bus_5c4dede9_;
input	[15:0]	bus_253147b9_;
input		bus_4ebaa98e_;
input	[15:0]	bus_5ceaaebb_;
input		bus_63833c02_;
input	[15:0]	bus_50790775_;
input		bus_2264995f_;
input	[15:0]	bus_1cdbfe01_;
input		bus_2c539ca8_;
input	[15:0]	bus_632c90cd_;
input		bus_2397b779_;
input	[15:0]	bus_26b5b1f6_;
input		bus_2570bc16_;
input	[15:0]	bus_48005bbe_;
input		bus_441deb71_;
input	[15:0]	bus_46b2645c_;
input		bus_62a23944_;
input	[15:0]	bus_1378e939_;
input		bus_513697cc_;
input	[15:0]	bus_2cee4380_;
input		bus_0475cc13_;
input	[15:0]	bus_78940204_;
input		bus_766fd037_;
input	[15:0]	bus_4d505dca_;
input		bus_1de90dae_;
input	[15:0]	bus_20ace7e3_;
input		bus_1c515fcc_;
input	[15:0]	bus_5e13118c_;
input		bus_041f2681_;
input	[15:0]	bus_6056c028_;
input		bus_3aa04241_;
input	[15:0]	bus_3321cb07_;
input		bus_7e50ec6c_;
input	[15:0]	bus_26d18263_;
output	[15:0]	bus_2a7d4abb_;
wire	[15:0]	endianswapper_077bd2d3_out;
wire		or_7bfb4760_u0;
wire	[15:0]	endianswapper_6f898fe2_out;
LL1_H_iunzipFilter2D_endianswapper_077bd2d3_ LL1_H_iunzipFilter2D_endianswapper_077bd2d3__1(.endianswapper_077bd2d3_in(16'h0), 
  .endianswapper_077bd2d3_out(endianswapper_077bd2d3_out));
assign bus_2a7d4abb_=16'h0;
assign or_7bfb4760_u0=bus_674bf37e_|bus_4a2d20e1_|bus_5c4dede9_|bus_4ebaa98e_|bus_63833c02_|bus_2264995f_|bus_2c539ca8_|bus_2397b779_|bus_2570bc16_|bus_441deb71_|bus_62a23944_|bus_513697cc_|bus_0475cc13_|bus_766fd037_|bus_1de90dae_|bus_1c515fcc_|bus_041f2681_|bus_3aa04241_|bus_7e50ec6c_;
LL1_H_iunzipFilter2D_endianswapper_6f898fe2_ LL1_H_iunzipFilter2D_endianswapper_6f898fe2__1(.endianswapper_6f898fe2_in(16'h0), 
  .endianswapper_6f898fe2_out(endianswapper_6f898fe2_out));
endmodule



module LL1_H_iunzipFilter2D_midRight2(CLK, RESET, GO, port_5ef6bce8_, port_5d219e2c_, port_7888f833_, port_0faf4797_, port_46e25d42_, port_5cd1a04c_, port_06fd2eaf_, RESULT, RESULT_u236, RESULT_u237, RESULT_u238, RESULT_u239, RESULT_u240, RESULT_u241, RESULT_u242, RESULT_u243, RESULT_u244, RESULT_u245, RESULT_u246, RESULT_u247, RESULT_u248, RESULT_u249, RESULT_u250, RESULT_u251, RESULT_u252, RESULT_u253, RESULT_u254, RESULT_u255, DONE);
input		CLK;
input		RESET;
input		GO;
input	[31:0]	port_5ef6bce8_;
input	[15:0]	port_5d219e2c_;
input		port_7888f833_;
input		port_0faf4797_;
input	[15:0]	port_46e25d42_;
input		port_5cd1a04c_;
input	[15:0]	port_06fd2eaf_;
output		RESULT;
output	[15:0]	RESULT_u236;
output		RESULT_u237;
output	[31:0]	RESULT_u238;
output		RESULT_u239;
output	[15:0]	RESULT_u240;
output		RESULT_u241;
output	[15:0]	RESULT_u242;
output		RESULT_u243;
output		RESULT_u244;
output		RESULT_u245;
output	[31:0]	RESULT_u246;
output	[2:0]	RESULT_u247;
output		RESULT_u248;
output	[31:0]	RESULT_u249;
output	[15:0]	RESULT_u250;
output	[2:0]	RESULT_u251;
output		RESULT_u252;
output	[15:0]	RESULT_u253;
output		RESULT_u254;
output	[15:0]	RESULT_u255;
output		DONE;
wire		simplePinWrite;
reg		done_cache_u28=1'h0;
wire		and_u312_u0;
wire		or_u67_u0;
wire		and_u317_u0;
wire		or_u68_u0;
reg		done_cache_u29_u0=1'h0;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_6ea17d98_instance_RESULT;
wire		or_u69_u0;
reg		reg_68249367_u0=1'h0;
wire		and_u326_u0;
wire	[31:0]	add;
wire	[15:0]	add_u6;
wire		not_u48;
wire		simplePinWrite_u61;
wire	[15:0]	simplePinWrite_u62;
wire	[15:0]	simplePinWrite_u63;
reg	[15:0]	syncEnable_u20=16'h0;
reg		reg_48151439_u0=1'h0;
reg		reg_48151439_result_delayed_u0=1'h0;
wire		or_u70_u0;
reg		reg_1be67ce5_u0=1'h0;
reg		reg_1817a137_u0=1'h0;
reg		reg_48151439_result_delayed_result_delayed_u0=1'h0;
reg	[15:0]	syncEnable_u21_u0=16'h0;
reg		reg_48151439_result_delayed_result_delayed_result_delayed_u0=1'h0;
assign simplePinWrite=GO&{1{GO}};
always @(posedge CLK or posedge GO or posedge or_u67_u0)
begin
if (or_u67_u0)
done_cache_u28<=1'h0;
else if (GO)
done_cache_u28<=1'h1;
else done_cache_u28<=done_cache_u28;
end
assign and_u312_u0=done_cache_u28&port_5cd1a04c_;
assign or_u67_u0=and_u312_u0|RESET;
assign and_u317_u0=done_cache_u29_u0&port_5cd1a04c_;
assign or_u68_u0=and_u317_u0|RESET;
always @(posedge CLK or posedge reg_1be67ce5_u0 or posedge or_u68_u0)
begin
if (or_u68_u0)
done_cache_u29_u0<=1'h0;
else if (reg_1be67ce5_u0)
done_cache_u29_u0<=1'h1;
else done_cache_u29_u0<=done_cache_u29_u0;
end
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_6ea17d98_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_6ea17d98_instance(.GO(reg_48151439_u0), 
  .port_7b5a94cd_(syncEnable_u20), .port_662c4c53_(port_46e25d42_), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_6ea17d98_instance_RESULT));
assign or_u69_u0=and_u326_u0|RESET;
always @(posedge CLK or posedge reg_48151439_result_delayed_result_delayed_u0 or posedge or_u69_u0)
begin
if (or_u69_u0)
reg_68249367_u0<=1'h0;
else if (reg_48151439_result_delayed_result_delayed_u0)
reg_68249367_u0<=1'h1;
else reg_68249367_u0<=reg_68249367_u0;
end
assign and_u326_u0=reg_68249367_u0&port_5cd1a04c_;
assign add=port_5ef6bce8_+32'h1;
assign add_u6=port_5d219e2c_+16'h1;
assign not_u48=!port_7888f833_;
assign simplePinWrite_u61=reg_48151439_u0&{1{reg_48151439_u0}};
assign simplePinWrite_u62=16'h1&{16{1'h1}};
assign simplePinWrite_u63=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_6ea17d98_instance_RESULT&{16{reg_48151439_u0}};
always @(posedge CLK)
begin
if (reg_1817a137_u0)
syncEnable_u20<=port_46e25d42_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_48151439_u0<=1'h0;
else reg_48151439_u0<=reg_1be67ce5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_48151439_result_delayed_u0<=1'h0;
else reg_48151439_result_delayed_u0<=reg_48151439_u0;
end
assign or_u70_u0=GO|reg_1be67ce5_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1be67ce5_u0<=1'h0;
else reg_1be67ce5_u0<=reg_1817a137_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1817a137_u0<=1'h0;
else reg_1817a137_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_48151439_result_delayed_result_delayed_u0<=1'h0;
else reg_48151439_result_delayed_result_delayed_u0<=reg_48151439_result_delayed_u0;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u21_u0<=port_06fd2eaf_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_48151439_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_48151439_result_delayed_result_delayed_result_delayed_u0<=reg_48151439_result_delayed_result_delayed_u0;
end
assign RESULT=GO;
assign RESULT_u236=16'h0;
assign RESULT_u237=GO;
assign RESULT_u238=add;
assign RESULT_u239=GO;
assign RESULT_u240=add_u6;
assign RESULT_u241=GO;
assign RESULT_u242=16'h0;
assign RESULT_u243=GO;
assign RESULT_u244=not_u48;
assign RESULT_u245=or_u70_u0;
assign RESULT_u246=32'h0;
assign RESULT_u247=3'h1;
assign RESULT_u248=reg_48151439_result_delayed_result_delayed_u0;
assign RESULT_u249=32'h0;
assign RESULT_u250=syncEnable_u21_u0;
assign RESULT_u251=3'h1;
assign RESULT_u252=simplePinWrite;
assign RESULT_u253=simplePinWrite_u62;
assign RESULT_u254=simplePinWrite_u61;
assign RESULT_u255=simplePinWrite_u63;
assign DONE=reg_48151439_result_delayed_result_delayed_result_delayed_u0;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_6ea17d98_(GO, port_7b5a94cd_, port_662c4c53_, RESULT);
input		GO;
input	[15:0]	port_7b5a94cd_;
input	[15:0]	port_662c4c53_;
output	[15:0]	RESULT;
wire	[15:0]	subtract;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_3792602a_instance_RESULT;
assign subtract=port_7b5a94cd_-port_662c4c53_;
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_3792602a_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_3792602a_instance(.GO(GO), 
  .port_17e78df6_({subtract[15], subtract[15:1]}), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_3792602a_instance_RESULT));
assign RESULT=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_3792602a_instance_RESULT;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_3792602a_(GO, port_17e78df6_, RESULT);
input		GO;
input	[15:0]	port_17e78df6_;
output	[15:0]	RESULT;
wire signed	[15:0]	greaterThan_a_signed;
wire signed	[15:0]	greaterThan_b_signed;
wire		greaterThan;
wire		and_u321_u0;
wire		and_u322_u0;
wire		not_u47_u0;
wire		and_u323_u0;
wire	[15:0]	mux_u23;
wire		and_u324_u0;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_17e78df6_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign and_u321_u0=GO&not_u47_u0;
assign and_u322_u0=GO&greaterThan;
assign not_u47_u0=~greaterThan;
assign and_u323_u0=and_u321_u0&GO;
assign mux_u23=(and_u323_u0)?port_17e78df6_:16'h0;
assign and_u324_u0=and_u322_u0&GO;
assign RESULT=mux_u23;
endmodule



module LL1_H_iunzipFilter2D_globalreset_physical_1f6e1ed4_(bus_68f6b794_, bus_1df2d7fb_, bus_23506230_);
input		bus_68f6b794_;
input		bus_1df2d7fb_;
output		bus_23506230_;
wire		or_2b5e0d8f_u0;
wire		and_7aff526d_u0;
wire		not_68e2b1d7_u0;
reg		sample_u6=1'h0;
reg		cross_u6=1'h0;
reg		glitch_u6=1'h0;
reg		final_u6=1'h1;
assign bus_23506230_=or_2b5e0d8f_u0;
assign or_2b5e0d8f_u0=bus_1df2d7fb_|final_u6;
assign and_7aff526d_u0=cross_u6&glitch_u6;
assign not_68e2b1d7_u0=~and_7aff526d_u0;
always @(posedge bus_68f6b794_)
begin
sample_u6<=1'h1;
end
always @(posedge bus_68f6b794_)
begin
cross_u6<=sample_u6;
end
always @(posedge bus_68f6b794_)
begin
glitch_u6<=cross_u6;
end
always @(posedge bus_68f6b794_)
begin
final_u6<=not_68e2b1d7_u0;
end
endmodule



module LL1_H_iunzipFilter2D_endianswapper_1ef5cadd_(endianswapper_1ef5cadd_in, endianswapper_1ef5cadd_out);
input	[15:0]	endianswapper_1ef5cadd_in;
output	[15:0]	endianswapper_1ef5cadd_out;
assign endianswapper_1ef5cadd_out=endianswapper_1ef5cadd_in;
endmodule



module LL1_H_iunzipFilter2D_endianswapper_5383acf9_(endianswapper_5383acf9_in, endianswapper_5383acf9_out);
input	[15:0]	endianswapper_5383acf9_in;
output	[15:0]	endianswapper_5383acf9_out;
assign endianswapper_5383acf9_out=endianswapper_5383acf9_in;
endmodule



module LL1_H_iunzipFilter2D_stateVar_processedRows(bus_50bd0603_, bus_06976a41_, bus_334b47c1_, bus_360674e9_, bus_2a00d576_, bus_52b2c6ce_, bus_5ab10369_, bus_7b0dad4e_, bus_691edc7e_, bus_2c378729_, bus_39e8dab6_, bus_22ec21fb_, bus_2bab2c65_, bus_4dee9c66_, bus_20abe20d_, bus_6396d044_, bus_47b99ec4_, bus_5b45ada7_, bus_4cb9b263_);
input		bus_50bd0603_;
input		bus_06976a41_;
input		bus_334b47c1_;
input	[15:0]	bus_360674e9_;
input		bus_2a00d576_;
input	[15:0]	bus_52b2c6ce_;
input		bus_5ab10369_;
input	[15:0]	bus_7b0dad4e_;
input		bus_691edc7e_;
input	[15:0]	bus_2c378729_;
input		bus_39e8dab6_;
input	[15:0]	bus_22ec21fb_;
input		bus_2bab2c65_;
input	[15:0]	bus_4dee9c66_;
input		bus_20abe20d_;
input	[15:0]	bus_6396d044_;
input		bus_47b99ec4_;
input	[15:0]	bus_5b45ada7_;
output	[15:0]	bus_4cb9b263_;
wire	[15:0]	mux_4019587a_u0;
wire		or_57d79e40_u0;
reg	[15:0]	stateVar_processedRows_u0=16'h0;
wire	[15:0]	endianswapper_1ef5cadd_out;
wire	[15:0]	endianswapper_5383acf9_out;
assign mux_4019587a_u0=({16{bus_334b47c1_}}&bus_360674e9_)|({16{bus_2a00d576_}}&16'h1)|({16{bus_5ab10369_}}&bus_7b0dad4e_)|({16{bus_691edc7e_}}&bus_2c378729_)|({16{bus_39e8dab6_}}&bus_22ec21fb_)|({16{bus_2bab2c65_}}&bus_4dee9c66_)|({16{bus_20abe20d_}}&16'h0)|({16{bus_47b99ec4_}}&16'h0);
assign bus_4cb9b263_=endianswapper_1ef5cadd_out;
assign or_57d79e40_u0=bus_334b47c1_|bus_2a00d576_|bus_5ab10369_|bus_691edc7e_|bus_39e8dab6_|bus_2bab2c65_|bus_20abe20d_|bus_47b99ec4_;
always @(posedge bus_50bd0603_ or posedge bus_06976a41_)
begin
if (bus_06976a41_)
stateVar_processedRows_u0<=16'h0;
else if (or_57d79e40_u0)
stateVar_processedRows_u0<=endianswapper_5383acf9_out;
end
LL1_H_iunzipFilter2D_endianswapper_1ef5cadd_ LL1_H_iunzipFilter2D_endianswapper_1ef5cadd__1(.endianswapper_1ef5cadd_in(stateVar_processedRows_u0), 
  .endianswapper_1ef5cadd_out(endianswapper_1ef5cadd_out));
LL1_H_iunzipFilter2D_endianswapper_5383acf9_ LL1_H_iunzipFilter2D_endianswapper_5383acf9__1(.endianswapper_5383acf9_in(mux_4019587a_u0), 
  .endianswapper_5383acf9_out(endianswapper_5383acf9_out));
endmodule



module LL1_H_iunzipFilter2D_bottomRightNoConsume2(CLK, RESET, GO, port_1379735b_, port_718e624c_, port_680823aa_, RESULT, RESULT_u256, RESULT_u257, RESULT_u258, RESULT_u259, RESULT_u260, RESULT_u261, RESULT_u262, RESULT_u263, RESULT_u264, RESULT_u265, RESULT_u266, RESULT_u267, RESULT_u268, RESULT_u269, RESULT_u270, DONE);
input		CLK;
input		RESET;
input		GO;
input		port_1379735b_;
input		port_718e624c_;
input	[15:0]	port_680823aa_;
output		RESULT;
output	[15:0]	RESULT_u256;
output		RESULT_u257;
output	[15:0]	RESULT_u258;
output		RESULT_u259;
output	[15:0]	RESULT_u260;
output		RESULT_u261;
output	[31:0]	RESULT_u262;
output		RESULT_u263;
output		RESULT_u264;
output		RESULT_u265;
output	[31:0]	RESULT_u266;
output	[2:0]	RESULT_u267;
output	[15:0]	RESULT_u268;
output		RESULT_u269;
output	[15:0]	RESULT_u270;
output		DONE;
reg		done_cache_u30=1'h0;
wire		and_u329_u0;
wire		or_u71_u0;
wire		and_u334_u0;
wire		or_u72_u0;
reg		done_cache_u31_u0=1'h0;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_04af7570_instance_RESULT;
wire		not_u50;
wire		simplePinWrite;
wire	[15:0]	simplePinWrite_u64;
wire	[15:0]	simplePinWrite_u65;
reg		reg_253c231b_u0=1'h0;
reg		reg_3e94c1ec_u0=1'h0;
reg		reg_47c9bc44_u0=1'h0;
reg		reg_3e94c1ec_result_delayed_u0=1'h0;
reg	[15:0]	syncEnable_u22=16'h0;
reg		reg_253c231b_result_delayed_u0=1'h0;
wire		or_u73_u0;
always @(posedge CLK or posedge GO or posedge or_u71_u0)
begin
if (or_u71_u0)
done_cache_u30<=1'h0;
else if (GO)
done_cache_u30<=1'h1;
else done_cache_u30<=done_cache_u30;
end
assign and_u329_u0=done_cache_u30&port_718e624c_;
assign or_u71_u0=and_u329_u0|RESET;
assign and_u334_u0=done_cache_u31_u0&port_718e624c_;
assign or_u72_u0=and_u334_u0|RESET;
always @(posedge CLK or posedge reg_253c231b_u0 or posedge or_u72_u0)
begin
if (or_u72_u0)
done_cache_u31_u0<=1'h0;
else if (reg_253c231b_u0)
done_cache_u31_u0<=1'h1;
else done_cache_u31_u0<=done_cache_u31_u0;
end
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_04af7570_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_04af7570_instance(.GO(reg_253c231b_result_delayed_u0), 
  .port_400ae17f_(syncEnable_u22), .port_14654d97_(port_680823aa_), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_04af7570_instance_RESULT));
assign not_u50=!port_1379735b_;
assign simplePinWrite=reg_253c231b_result_delayed_u0&{1{reg_253c231b_result_delayed_u0}};
assign simplePinWrite_u64=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_04af7570_instance_RESULT&{16{reg_253c231b_result_delayed_u0}};
assign simplePinWrite_u65=16'h1&{16{1'h1}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_253c231b_u0<=1'h0;
else reg_253c231b_u0<=reg_47c9bc44_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3e94c1ec_u0<=1'h0;
else reg_3e94c1ec_u0<=reg_253c231b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_47c9bc44_u0<=1'h0;
else reg_47c9bc44_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3e94c1ec_result_delayed_u0<=1'h0;
else reg_3e94c1ec_result_delayed_u0<=reg_3e94c1ec_u0;
end
always @(posedge CLK)
begin
if (reg_47c9bc44_u0)
syncEnable_u22<=port_680823aa_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_253c231b_result_delayed_u0<=1'h0;
else reg_253c231b_result_delayed_u0<=reg_253c231b_u0;
end
assign or_u73_u0=GO|reg_253c231b_u0;
assign RESULT=GO;
assign RESULT_u256=16'h0;
assign RESULT_u257=GO;
assign RESULT_u258=16'h0;
assign RESULT_u259=GO;
assign RESULT_u260=16'h0;
assign RESULT_u261=GO;
assign RESULT_u262=32'h0;
assign RESULT_u263=GO;
assign RESULT_u264=not_u50;
assign RESULT_u265=or_u73_u0;
assign RESULT_u266=32'h0;
assign RESULT_u267=3'h1;
assign RESULT_u268=simplePinWrite_u65;
assign RESULT_u269=simplePinWrite;
assign RESULT_u270=simplePinWrite_u64;
assign DONE=reg_3e94c1ec_result_delayed_u0;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_04af7570_(GO, port_400ae17f_, port_14654d97_, RESULT);
input		GO;
input	[15:0]	port_400ae17f_;
input	[15:0]	port_14654d97_;
output	[15:0]	RESULT;
wire	[15:0]	subtract;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_6e000804_instance_RESULT;
assign subtract=port_400ae17f_-port_14654d97_;
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_6e000804_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_6e000804_instance(.GO(GO), 
  .port_08fc5cfc_({subtract[15], subtract[15:1]}), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_6e000804_instance_RESULT));
assign RESULT=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_6e000804_instance_RESULT;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_6e000804_(GO, port_08fc5cfc_, RESULT);
input		GO;
input	[15:0]	port_08fc5cfc_;
output	[15:0]	RESULT;
wire signed	[15:0]	greaterThan_b_signed;
wire		greaterThan;
wire signed	[15:0]	greaterThan_a_signed;
wire		and_u338_u0;
wire		not_u49_u0;
wire		and_u339_u0;
wire		and_u340_u0;
wire	[15:0]	mux_u24;
wire		and_u341_u0;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_08fc5cfc_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign and_u338_u0=GO&greaterThan;
assign not_u49_u0=~greaterThan;
assign and_u339_u0=GO&not_u49_u0;
assign and_u340_u0=and_u339_u0&GO;
assign mux_u24=(and_u341_u0)?16'h0:port_08fc5cfc_;
assign and_u341_u0=and_u338_u0&GO;
assign RESULT=mux_u24;
endmodule



module LL1_H_iunzipFilter2D_mid2(CLK, RESET, GO, port_63ca52d3_, port_3ed342e9_, port_61009e2d_, port_5174b1c2_, port_22e17dd6_, port_28805c0d_, RESULT, RESULT_u271, RESULT_u272, RESULT_u273, RESULT_u274, RESULT_u275, RESULT_u276, RESULT_u277, RESULT_u278, RESULT_u279, RESULT_u280, RESULT_u281, RESULT_u282, RESULT_u283, RESULT_u284, RESULT_u285, RESULT_u286, DONE);
input		CLK;
input		RESET;
input		GO;
input	[31:0]	port_63ca52d3_;
input	[15:0]	port_3ed342e9_;
input		port_61009e2d_;
input	[15:0]	port_5174b1c2_;
input		port_22e17dd6_;
input	[15:0]	port_28805c0d_;
output		RESULT;
output	[31:0]	RESULT_u271;
output		RESULT_u272;
output	[15:0]	RESULT_u273;
output		RESULT_u274;
output	[15:0]	RESULT_u275;
output		RESULT_u276;
output	[31:0]	RESULT_u277;
output	[2:0]	RESULT_u278;
output		RESULT_u279;
output	[31:0]	RESULT_u280;
output	[15:0]	RESULT_u281;
output	[2:0]	RESULT_u282;
output		RESULT_u283;
output	[15:0]	RESULT_u284;
output	[15:0]	RESULT_u285;
output		RESULT_u286;
output		DONE;
wire		simplePinWrite;
reg		done_cache_u32=1'h0;
wire		or_u74_u0;
wire		and_u343_u0;
wire		and_u348_u0;
wire		or_u75_u0;
reg		done_cache_u33_u0=1'h0;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_5ef1d326_instance_RESULT;
wire		or_u76_u0;
reg		reg_213565e9_u0=1'h0;
wire		and_u357_u0;
wire	[31:0]	add;
wire	[15:0]	add_u7;
wire	[15:0]	simplePinWrite_u66;
wire	[15:0]	simplePinWrite_u67;
wire		simplePinWrite_u68;
reg	[15:0]	syncEnable_u23=16'h0;
reg		reg_065194d2_u0=1'h0;
wire		or_u77_u0;
reg		reg_664b6a80_u0=1'h0;
reg	[15:0]	syncEnable_u24_u0=16'h0;
reg		reg_6a7bff7c_u0=1'h0;
reg		reg_065194d2_result_delayed_u0=1'h0;
reg		reg_664b6a80_result_delayed_u0=1'h0;
reg		reg_664b6a80_result_delayed_result_delayed_u0=1'h0;
assign simplePinWrite=GO&{1{GO}};
always @(posedge CLK or posedge GO or posedge or_u74_u0)
begin
if (or_u74_u0)
done_cache_u32<=1'h0;
else if (GO)
done_cache_u32<=1'h1;
else done_cache_u32<=done_cache_u32;
end
assign or_u74_u0=and_u343_u0|RESET;
assign and_u343_u0=done_cache_u32&port_22e17dd6_;
assign and_u348_u0=done_cache_u33_u0&port_22e17dd6_;
assign or_u75_u0=and_u348_u0|RESET;
always @(posedge CLK or posedge reg_065194d2_u0 or posedge or_u75_u0)
begin
if (or_u75_u0)
done_cache_u33_u0<=1'h0;
else if (reg_065194d2_u0)
done_cache_u33_u0<=1'h1;
else done_cache_u33_u0<=done_cache_u33_u0;
end
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_5ef1d326_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_5ef1d326_instance(.GO(reg_065194d2_result_delayed_u0), 
  .port_6aa520ec_(syncEnable_u24_u0), .port_3f5c5b34_(port_5174b1c2_), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_5ef1d326_instance_RESULT));
assign or_u76_u0=and_u357_u0|RESET;
always @(posedge CLK or posedge reg_664b6a80_result_delayed_u0 or posedge or_u76_u0)
begin
if (or_u76_u0)
reg_213565e9_u0<=1'h0;
else if (reg_664b6a80_result_delayed_u0)
reg_213565e9_u0<=1'h1;
else reg_213565e9_u0<=reg_213565e9_u0;
end
assign and_u357_u0=reg_213565e9_u0&port_22e17dd6_;
assign add=port_63ca52d3_+32'h1;
assign add_u7=port_3ed342e9_+16'h1;
assign simplePinWrite_u66=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_5ef1d326_instance_RESULT&{16{reg_065194d2_result_delayed_u0}};
assign simplePinWrite_u67=16'h1&{16{1'h1}};
assign simplePinWrite_u68=reg_065194d2_result_delayed_u0&{1{reg_065194d2_result_delayed_u0}};
always @(posedge CLK)
begin
if (GO)
syncEnable_u23<=port_28805c0d_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_065194d2_u0<=1'h0;
else reg_065194d2_u0<=reg_6a7bff7c_u0;
end
assign or_u77_u0=GO|reg_065194d2_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_664b6a80_u0<=1'h0;
else reg_664b6a80_u0<=reg_065194d2_result_delayed_u0;
end
always @(posedge CLK)
begin
if (reg_6a7bff7c_u0)
syncEnable_u24_u0<=port_5174b1c2_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6a7bff7c_u0<=1'h0;
else reg_6a7bff7c_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_065194d2_result_delayed_u0<=1'h0;
else reg_065194d2_result_delayed_u0<=reg_065194d2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_664b6a80_result_delayed_u0<=1'h0;
else reg_664b6a80_result_delayed_u0<=reg_664b6a80_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_664b6a80_result_delayed_result_delayed_u0<=1'h0;
else reg_664b6a80_result_delayed_result_delayed_u0<=reg_664b6a80_result_delayed_u0;
end
assign RESULT=GO;
assign RESULT_u271=add;
assign RESULT_u272=GO;
assign RESULT_u273=16'h0;
assign RESULT_u274=GO;
assign RESULT_u275=add_u7;
assign RESULT_u276=or_u77_u0;
assign RESULT_u277=32'h0;
assign RESULT_u278=3'h1;
assign RESULT_u279=reg_664b6a80_result_delayed_u0;
assign RESULT_u280=32'h0;
assign RESULT_u281=syncEnable_u23;
assign RESULT_u282=3'h1;
assign RESULT_u283=simplePinWrite;
assign RESULT_u284=simplePinWrite_u67;
assign RESULT_u285=simplePinWrite_u66;
assign RESULT_u286=simplePinWrite_u68;
assign DONE=reg_664b6a80_result_delayed_result_delayed_u0;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_5ef1d326_(GO, port_6aa520ec_, port_3f5c5b34_, RESULT);
input		GO;
input	[15:0]	port_6aa520ec_;
input	[15:0]	port_3f5c5b34_;
output	[15:0]	RESULT;
wire	[15:0]	subtract;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_65475dd0_instance_RESULT;
assign subtract=port_6aa520ec_-port_3f5c5b34_;
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_65475dd0_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_65475dd0_instance(.GO(GO), 
  .port_18babcf0_({subtract[15], subtract[15:1]}), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_65475dd0_instance_RESULT));
assign RESULT=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_65475dd0_instance_RESULT;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_65475dd0_(GO, port_18babcf0_, RESULT);
input		GO;
input	[15:0]	port_18babcf0_;
output	[15:0]	RESULT;
wire		greaterThan;
wire signed	[15:0]	greaterThan_b_signed;
wire signed	[15:0]	greaterThan_a_signed;
wire		not_u51_u0;
wire		and_u352_u0;
wire		and_u353_u0;
wire		and_u354_u0;
wire	[15:0]	mux_u25;
wire		and_u355_u0;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_18babcf0_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign not_u51_u0=~greaterThan;
assign and_u352_u0=GO&not_u51_u0;
assign and_u353_u0=GO&greaterThan;
assign and_u354_u0=and_u353_u0&GO;
assign mux_u25=(and_u354_u0)?16'h0:port_18babcf0_;
assign and_u355_u0=and_u352_u0&GO;
assign RESULT=mux_u25;
endmodule



module LL1_H_iunzipFilter2D_bottomRowNoConsume2(CLK, RESET, GO, port_0c13a378_, port_55afd2df_, port_137c836d_, RESULT, RESULT_u287, RESULT_u288, RESULT_u289, RESULT_u290, RESULT_u291, RESULT_u292, RESULT_u293, RESULT_u294, RESULT_u295, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_0c13a378_;
input		port_55afd2df_;
input	[15:0]	port_137c836d_;
output		RESULT;
output	[15:0]	RESULT_u287;
output		RESULT_u288;
output	[15:0]	RESULT_u289;
output		RESULT_u290;
output	[31:0]	RESULT_u291;
output	[2:0]	RESULT_u292;
output	[15:0]	RESULT_u293;
output	[15:0]	RESULT_u294;
output		RESULT_u295;
output		DONE;
reg		done_cache_u34=1'h0;
wire		and_u360_u0;
wire		or_u78_u0;
wire		and_u365_u0;
reg		done_cache_u35_u0=1'h0;
wire		or_u79_u0;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_58c8fd93_instance_RESULT;
wire	[15:0]	add;
wire	[15:0]	simplePinWrite;
wire	[15:0]	simplePinWrite_u69;
wire		simplePinWrite_u70;
reg		reg_73979caf_u0=1'h0;
reg		reg_722de161_u0=1'h0;
wire		or_u80_u0;
reg	[15:0]	syncEnable_u25=16'h0;
reg		reg_5882f729_u0=1'h0;
reg		reg_722de161_result_delayed_u0=1'h0;
reg		reg_73979caf_result_delayed_u0=1'h0;
always @(posedge CLK or posedge GO or posedge or_u78_u0)
begin
if (or_u78_u0)
done_cache_u34<=1'h0;
else if (GO)
done_cache_u34<=1'h1;
else done_cache_u34<=done_cache_u34;
end
assign and_u360_u0=done_cache_u34&port_55afd2df_;
assign or_u78_u0=and_u360_u0|RESET;
assign and_u365_u0=done_cache_u35_u0&port_55afd2df_;
always @(posedge CLK or posedge reg_73979caf_result_delayed_u0 or posedge or_u79_u0)
begin
if (or_u79_u0)
done_cache_u35_u0<=1'h0;
else if (reg_73979caf_result_delayed_u0)
done_cache_u35_u0<=1'h1;
else done_cache_u35_u0<=done_cache_u35_u0;
end
assign or_u79_u0=and_u365_u0|RESET;
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_58c8fd93_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_58c8fd93_instance(.GO(reg_5882f729_u0), 
  .port_009aaf7b_(syncEnable_u25), .port_10414408_(port_137c836d_), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_58c8fd93_instance_RESULT));
assign add=port_0c13a378_+16'h1;
assign simplePinWrite=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_58c8fd93_instance_RESULT&{16{reg_5882f729_u0}};
assign simplePinWrite_u69=16'h1&{16{1'h1}};
assign simplePinWrite_u70=reg_5882f729_u0&{1{reg_5882f729_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_73979caf_u0<=1'h0;
else reg_73979caf_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_722de161_u0<=1'h0;
else reg_722de161_u0<=reg_5882f729_u0;
end
assign or_u80_u0=GO|reg_73979caf_result_delayed_u0;
always @(posedge CLK)
begin
if (reg_73979caf_u0)
syncEnable_u25<=port_137c836d_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5882f729_u0<=1'h0;
else reg_5882f729_u0<=reg_73979caf_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_722de161_result_delayed_u0<=1'h0;
else reg_722de161_result_delayed_u0<=reg_722de161_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_73979caf_result_delayed_u0<=1'h0;
else reg_73979caf_result_delayed_u0<=reg_73979caf_u0;
end
assign RESULT=GO;
assign RESULT_u287=16'h0;
assign RESULT_u288=GO;
assign RESULT_u289=add;
assign RESULT_u290=or_u80_u0;
assign RESULT_u291=32'h0;
assign RESULT_u292=3'h1;
assign RESULT_u293=simplePinWrite_u69;
assign RESULT_u294=simplePinWrite;
assign RESULT_u295=simplePinWrite_u70;
assign DONE=reg_722de161_result_delayed_u0;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_58c8fd93_(GO, port_009aaf7b_, port_10414408_, RESULT);
input		GO;
input	[15:0]	port_009aaf7b_;
input	[15:0]	port_10414408_;
output	[15:0]	RESULT;
wire	[15:0]	subtract;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_2b524786_instance_RESULT;
assign subtract=port_009aaf7b_-port_10414408_;
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_2b524786_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_2b524786_instance(.GO(GO), 
  .port_0a50b3b6_({subtract[15], subtract[15:1]}), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_2b524786_instance_RESULT));
assign RESULT=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_2b524786_instance_RESULT;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_2b524786_(GO, port_0a50b3b6_, RESULT);
input		GO;
input	[15:0]	port_0a50b3b6_;
output	[15:0]	RESULT;
wire signed	[15:0]	greaterThan_a_signed;
wire		greaterThan;
wire signed	[15:0]	greaterThan_b_signed;
wire		and_u369_u0;
wire		and_u370_u0;
wire		not_u52_u0;
wire		and_u371_u0;
wire	[15:0]	mux_u26;
wire		and_u372_u0;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_0a50b3b6_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign and_u369_u0=GO&greaterThan;
assign and_u370_u0=GO&not_u52_u0;
assign not_u52_u0=~greaterThan;
assign and_u371_u0=and_u369_u0&GO;
assign mux_u26=(and_u372_u0)?port_0a50b3b6_:16'h0;
assign and_u372_u0=and_u370_u0&GO;
assign RESULT=mux_u26;
endmodule



module LL1_H_iunzipFilter2D_midLeft2(CLK, RESET, GO, port_55a161f7_, port_7ef80ea3_, port_0e0f96e7_, port_425dfc12_, port_1c2a9de3_, port_7b60df17_, port_17ab7fa3_, RESULT, RESULT_u296, RESULT_u297, RESULT_u298, RESULT_u299, RESULT_u300, RESULT_u301, RESULT_u302, RESULT_u303, RESULT_u304, RESULT_u305, RESULT_u306, RESULT_u307, RESULT_u308, RESULT_u309, RESULT_u310, RESULT_u311, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_55a161f7_;
input	[31:0]	port_7ef80ea3_;
input	[15:0]	port_0e0f96e7_;
input		port_425dfc12_;
input	[15:0]	port_1c2a9de3_;
input		port_7b60df17_;
input	[15:0]	port_17ab7fa3_;
output		RESULT;
output	[15:0]	RESULT_u296;
output		RESULT_u297;
output	[31:0]	RESULT_u298;
output		RESULT_u299;
output	[15:0]	RESULT_u300;
output		RESULT_u301;
output	[31:0]	RESULT_u302;
output	[2:0]	RESULT_u303;
output		RESULT_u304;
output	[31:0]	RESULT_u305;
output	[15:0]	RESULT_u306;
output	[2:0]	RESULT_u307;
output		RESULT_u308;
output	[15:0]	RESULT_u309;
output		RESULT_u310;
output	[15:0]	RESULT_u311;
output		DONE;
wire		simplePinWrite;
reg		done_cache_u36=1'h0;
wire		and_u374_u0;
wire		or_u81_u0;
wire		and_u379_u0;
wire		or_u82_u0;
reg		done_cache_u37_u0=1'h0;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_3c3b5e00_instance_RESULT;
wire		or_u83_u0;
reg		reg_52bb81ec_u0=1'h0;
wire		and_u388_u0;
wire	[31:0]	add;
wire	[15:0]	add_u8;
wire		simplePinWrite_u71;
wire	[15:0]	simplePinWrite_u72;
wire	[15:0]	simplePinWrite_u73;
reg	[15:0]	syncEnable_u26=16'h0;
wire		or_u84_u0;
reg		reg_5f9682d1_u0=1'h0;
reg	[15:0]	syncEnable_u27_u0=16'h0;
reg		reg_5cd8e16e_u0=1'h0;
reg		reg_37bd2061_u0=1'h0;
reg		reg_5cd8e16e_result_delayed_u0=1'h0;
reg		reg_5f9682d1_result_delayed_u0=1'h0;
reg		reg_5f9682d1_result_delayed_result_delayed_u0=1'h0;
assign simplePinWrite=GO&{1{GO}};
always @(posedge CLK or posedge GO or posedge or_u81_u0)
begin
if (or_u81_u0)
done_cache_u36<=1'h0;
else if (GO)
done_cache_u36<=1'h1;
else done_cache_u36<=done_cache_u36;
end
assign and_u374_u0=done_cache_u36&port_7b60df17_;
assign or_u81_u0=and_u374_u0|RESET;
assign and_u379_u0=done_cache_u37_u0&port_7b60df17_;
assign or_u82_u0=and_u379_u0|RESET;
always @(posedge CLK or posedge reg_5cd8e16e_result_delayed_u0 or posedge or_u82_u0)
begin
if (or_u82_u0)
done_cache_u37_u0<=1'h0;
else if (reg_5cd8e16e_result_delayed_u0)
done_cache_u37_u0<=1'h1;
else done_cache_u37_u0<=done_cache_u37_u0;
end
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_3c3b5e00_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_3c3b5e00_instance(.GO(reg_5f9682d1_u0), 
  .port_0c6e9a0d_(syncEnable_u26), .port_6b73e1b7_(port_1c2a9de3_), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_3c3b5e00_instance_RESULT));
assign or_u83_u0=and_u388_u0|RESET;
always @(posedge CLK or posedge reg_5f9682d1_result_delayed_result_delayed_u0 or posedge or_u83_u0)
begin
if (or_u83_u0)
reg_52bb81ec_u0<=1'h0;
else if (reg_5f9682d1_result_delayed_result_delayed_u0)
reg_52bb81ec_u0<=1'h1;
else reg_52bb81ec_u0<=reg_52bb81ec_u0;
end
assign and_u388_u0=reg_52bb81ec_u0&port_7b60df17_;
assign add=port_7ef80ea3_+32'h1;
assign add_u8=port_0e0f96e7_+16'h1;
assign simplePinWrite_u71=reg_5f9682d1_u0&{1{reg_5f9682d1_u0}};
assign simplePinWrite_u72=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_3c3b5e00_instance_RESULT&{16{reg_5f9682d1_u0}};
assign simplePinWrite_u73=16'h1&{16{1'h1}};
always @(posedge CLK)
begin
if (reg_5cd8e16e_u0)
syncEnable_u26<=port_1c2a9de3_;
end
assign or_u84_u0=GO|reg_5cd8e16e_result_delayed_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5f9682d1_u0<=1'h0;
else reg_5f9682d1_u0<=reg_5cd8e16e_result_delayed_u0;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u27_u0<=port_17ab7fa3_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5cd8e16e_u0<=1'h0;
else reg_5cd8e16e_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_37bd2061_u0<=1'h0;
else reg_37bd2061_u0<=reg_5f9682d1_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5cd8e16e_result_delayed_u0<=1'h0;
else reg_5cd8e16e_result_delayed_u0<=reg_5cd8e16e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5f9682d1_result_delayed_u0<=1'h0;
else reg_5f9682d1_result_delayed_u0<=reg_5f9682d1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5f9682d1_result_delayed_result_delayed_u0<=1'h0;
else reg_5f9682d1_result_delayed_result_delayed_u0<=reg_5f9682d1_result_delayed_u0;
end
assign RESULT=GO;
assign RESULT_u296=16'h0;
assign RESULT_u297=GO;
assign RESULT_u298=add;
assign RESULT_u299=GO;
assign RESULT_u300=add_u8;
assign RESULT_u301=or_u84_u0;
assign RESULT_u302=32'h0;
assign RESULT_u303=3'h1;
assign RESULT_u304=reg_5f9682d1_result_delayed_result_delayed_u0;
assign RESULT_u305=32'h0;
assign RESULT_u306=syncEnable_u27_u0;
assign RESULT_u307=3'h1;
assign RESULT_u308=simplePinWrite;
assign RESULT_u309=simplePinWrite_u73;
assign RESULT_u310=simplePinWrite_u71;
assign RESULT_u311=simplePinWrite_u72;
assign DONE=reg_37bd2061_u0;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_3c3b5e00_(GO, port_0c6e9a0d_, port_6b73e1b7_, RESULT);
input		GO;
input	[15:0]	port_0c6e9a0d_;
input	[15:0]	port_6b73e1b7_;
output	[15:0]	RESULT;
wire	[15:0]	subtract;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_5eaeabee_instance_RESULT;
assign subtract=port_0c6e9a0d_-port_6b73e1b7_;
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_5eaeabee_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_5eaeabee_instance(.GO(GO), 
  .port_4cdcdf75_({subtract[15], subtract[15:1]}), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_5eaeabee_instance_RESULT));
assign RESULT=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_5eaeabee_instance_RESULT;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_5eaeabee_(GO, port_4cdcdf75_, RESULT);
input		GO;
input	[15:0]	port_4cdcdf75_;
output	[15:0]	RESULT;
wire signed	[15:0]	greaterThan_a_signed;
wire		greaterThan;
wire signed	[15:0]	greaterThan_b_signed;
wire		and_u383_u0;
wire		not_u53_u0;
wire		and_u384_u0;
wire	[15:0]	mux_u27;
wire		and_u385_u0;
wire		and_u386_u0;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_4cdcdf75_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign and_u383_u0=GO&not_u53_u0;
assign not_u53_u0=~greaterThan;
assign and_u384_u0=GO&greaterThan;
assign mux_u27=(and_u386_u0)?port_4cdcdf75_:16'h0;
assign and_u385_u0=and_u384_u0&GO;
assign and_u386_u0=and_u383_u0&GO;
assign RESULT=mux_u27;
endmodule



module LL1_H_iunzipFilter2D_endianswapper_596173d3_(endianswapper_596173d3_in, endianswapper_596173d3_out);
input	[31:0]	endianswapper_596173d3_in;
output	[31:0]	endianswapper_596173d3_out;
assign endianswapper_596173d3_out=endianswapper_596173d3_in;
endmodule



module LL1_H_iunzipFilter2D_endianswapper_349f28e3_(endianswapper_349f28e3_in, endianswapper_349f28e3_out);
input	[31:0]	endianswapper_349f28e3_in;
output	[31:0]	endianswapper_349f28e3_out;
assign endianswapper_349f28e3_out=endianswapper_349f28e3_in;
endmodule



module LL1_H_iunzipFilter2D_stateVar_consumed(bus_29e3f084_, bus_3ddb8871_, bus_41726d12_, bus_16da44fd_, bus_742d05ab_, bus_594dfb2b_, bus_4c0950d8_, bus_4229c30d_, bus_3cf40804_, bus_1b391612_, bus_553e65f0_, bus_35213476_, bus_6df9cec0_, bus_6e3ac2bf_, bus_777f8403_, bus_3b684d2d_, bus_7ad94f9e_, bus_7a612d89_, bus_57752a3a_, bus_6f16944e_, bus_77ad45a1_, bus_7708085a_, bus_5f8514a9_, bus_7ee2b5b9_, bus_0da1a829_, bus_56da0d80_, bus_69808cf7_);
input		bus_29e3f084_;
input		bus_3ddb8871_;
input		bus_41726d12_;
input	[31:0]	bus_16da44fd_;
input		bus_742d05ab_;
input	[31:0]	bus_594dfb2b_;
input		bus_4c0950d8_;
input	[31:0]	bus_4229c30d_;
input		bus_3cf40804_;
input	[31:0]	bus_1b391612_;
input		bus_553e65f0_;
input	[31:0]	bus_35213476_;
input		bus_6df9cec0_;
input	[31:0]	bus_6e3ac2bf_;
input		bus_777f8403_;
input	[31:0]	bus_3b684d2d_;
input		bus_7ad94f9e_;
input	[31:0]	bus_7a612d89_;
input		bus_57752a3a_;
input	[31:0]	bus_6f16944e_;
input		bus_77ad45a1_;
input	[31:0]	bus_7708085a_;
input		bus_5f8514a9_;
input	[31:0]	bus_7ee2b5b9_;
input		bus_0da1a829_;
input	[31:0]	bus_56da0d80_;
output	[31:0]	bus_69808cf7_;
wire	[31:0]	endianswapper_596173d3_out;
wire	[31:0]	mux_73c75d2c_u0;
reg	[31:0]	stateVar_consumed_u0=32'h0;
wire	[31:0]	endianswapper_349f28e3_out;
wire		or_2000cf5d_u0;
LL1_H_iunzipFilter2D_endianswapper_596173d3_ LL1_H_iunzipFilter2D_endianswapper_596173d3__1(.endianswapper_596173d3_in(mux_73c75d2c_u0), 
  .endianswapper_596173d3_out(endianswapper_596173d3_out));
assign bus_69808cf7_=endianswapper_349f28e3_out;
assign mux_73c75d2c_u0=({32{bus_41726d12_}}&bus_16da44fd_)|({32{bus_742d05ab_}}&bus_594dfb2b_)|({32{bus_4c0950d8_}}&bus_4229c30d_)|({32{bus_3cf40804_}}&bus_1b391612_)|({32{bus_553e65f0_}}&bus_35213476_)|({32{bus_6df9cec0_}}&bus_6e3ac2bf_)|({32{bus_777f8403_}}&bus_3b684d2d_)|({32{bus_7ad94f9e_}}&bus_7a612d89_)|({32{bus_57752a3a_}}&bus_6f16944e_)|({32{bus_77ad45a1_}}&bus_7708085a_)|({32{bus_5f8514a9_}}&32'h0)|({32{bus_0da1a829_}}&32'h0);
always @(posedge bus_29e3f084_ or posedge bus_3ddb8871_)
begin
if (bus_3ddb8871_)
stateVar_consumed_u0<=32'h0;
else if (or_2000cf5d_u0)
stateVar_consumed_u0<=endianswapper_596173d3_out;
end
LL1_H_iunzipFilter2D_endianswapper_349f28e3_ LL1_H_iunzipFilter2D_endianswapper_349f28e3__1(.endianswapper_349f28e3_in(stateVar_consumed_u0), 
  .endianswapper_349f28e3_out(endianswapper_349f28e3_out));
assign or_2000cf5d_u0=bus_41726d12_|bus_742d05ab_|bus_4c0950d8_|bus_3cf40804_|bus_553e65f0_|bus_6df9cec0_|bus_777f8403_|bus_7ad94f9e_|bus_57752a3a_|bus_77ad45a1_|bus_5f8514a9_|bus_0da1a829_;
endmodule



module LL1_H_iunzipFilter2D_endianswapper_53578707_(endianswapper_53578707_in, endianswapper_53578707_out);
input	[15:0]	endianswapper_53578707_in;
output	[15:0]	endianswapper_53578707_out;
assign endianswapper_53578707_out=endianswapper_53578707_in;
endmodule



module LL1_H_iunzipFilter2D_endianswapper_3523ce26_(endianswapper_3523ce26_in, endianswapper_3523ce26_out);
input	[15:0]	endianswapper_3523ce26_in;
output	[15:0]	endianswapper_3523ce26_out;
assign endianswapper_3523ce26_out=endianswapper_3523ce26_in;
endmodule



module LL1_H_iunzipFilter2D_stateVar_populatePtr(bus_42988fd2_, bus_63643b3f_, bus_65cf25d9_, bus_21d0a234_, bus_5fdc3a92_, bus_668e6817_, bus_70eb3e5c_);
input		bus_42988fd2_;
input		bus_63643b3f_;
input		bus_65cf25d9_;
input	[15:0]	bus_21d0a234_;
input		bus_5fdc3a92_;
input	[15:0]	bus_668e6817_;
output	[15:0]	bus_70eb3e5c_;
wire	[15:0]	endianswapper_53578707_out;
reg	[15:0]	stateVar_populatePtr_u0=16'h0;
wire	[15:0]	endianswapper_3523ce26_out;
wire	[15:0]	mux_3049bb9e_u0;
wire		or_58bc3e37_u0;
LL1_H_iunzipFilter2D_endianswapper_53578707_ LL1_H_iunzipFilter2D_endianswapper_53578707__1(.endianswapper_53578707_in(mux_3049bb9e_u0), 
  .endianswapper_53578707_out(endianswapper_53578707_out));
always @(posedge bus_42988fd2_ or posedge bus_63643b3f_)
begin
if (bus_63643b3f_)
stateVar_populatePtr_u0<=16'h0;
else if (or_58bc3e37_u0)
stateVar_populatePtr_u0<=endianswapper_53578707_out;
end
LL1_H_iunzipFilter2D_endianswapper_3523ce26_ LL1_H_iunzipFilter2D_endianswapper_3523ce26__1(.endianswapper_3523ce26_in(stateVar_populatePtr_u0), 
  .endianswapper_3523ce26_out(endianswapper_3523ce26_out));
assign mux_3049bb9e_u0=(bus_65cf25d9_)?bus_21d0a234_:16'h0;
assign bus_70eb3e5c_=endianswapper_3523ce26_out;
assign or_58bc3e37_u0=bus_65cf25d9_|bus_5fdc3a92_;
endmodule



module LL1_H_iunzipFilter2D_populateBuffer(CLK, RESET, GO, port_623c9ece_, port_165a8581_, port_7b608cd9_, port_4da138d8_, RESULT, RESULT_u312, RESULT_u313, RESULT_u314, RESULT_u315, RESULT_u316, RESULT_u317, RESULT_u318, RESULT_u319, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_623c9ece_;
input	[31:0]	port_165a8581_;
input		port_7b608cd9_;
input	[15:0]	port_4da138d8_;
output		RESULT;
output	[15:0]	RESULT_u312;
output		RESULT_u313;
output	[31:0]	RESULT_u314;
output		RESULT_u315;
output	[31:0]	RESULT_u316;
output	[15:0]	RESULT_u317;
output	[2:0]	RESULT_u318;
output		RESULT_u319;
output		DONE;
wire		simplePinWrite;
wire	[31:0]	add;
wire		and_u390_u0;
wire		or_u85_u0;
reg		reg_6c28de12_u0=1'h0;
wire	[31:0]	add_u9;
wire	[15:0]	add_u10;
reg		reg_479ac81b_u0=1'h0;
assign simplePinWrite=GO&{1{GO}};
assign add={port_623c9ece_[15], port_623c9ece_[15], port_623c9ece_[15], port_623c9ece_[15], port_623c9ece_[15], port_623c9ece_[15], port_623c9ece_[15], port_623c9ece_[15], port_623c9ece_[15], port_623c9ece_[15], port_623c9ece_[15], port_623c9ece_[15], port_623c9ece_[15], port_623c9ece_[15], port_623c9ece_[15], port_623c9ece_[15], port_623c9ece_}+32'h0;
assign and_u390_u0=reg_6c28de12_u0&port_7b608cd9_;
assign or_u85_u0=and_u390_u0|RESET;
always @(posedge CLK or posedge GO or posedge or_u85_u0)
begin
if (or_u85_u0)
reg_6c28de12_u0<=1'h0;
else if (GO)
reg_6c28de12_u0<=1'h1;
else reg_6c28de12_u0<=reg_6c28de12_u0;
end
assign add_u9=port_165a8581_+32'h1;
assign add_u10=port_623c9ece_+16'h1;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_479ac81b_u0<=1'h0;
else reg_479ac81b_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u312=add_u10;
assign RESULT_u313=GO;
assign RESULT_u314=add_u9;
assign RESULT_u315=GO;
assign RESULT_u316=add;
assign RESULT_u317=port_4da138d8_;
assign RESULT_u318=3'h1;
assign RESULT_u319=simplePinWrite;
assign DONE=reg_479ac81b_u0;
endmodule



module LL1_H_iunzipFilter2D_scheduler(CLK, RESET, GO, port_42620ba7_, port_41492b7c_, port_34f62b85_, port_6d2bfa2d_, port_2e0d86cd_, port_70e1f405_, port_6d3af1f9_, port_459c8efa_, port_24157214_, port_6e290ca0_, port_28187583_, port_5cc4abf1_, port_010adde4_, port_756b4eaa_, port_6004d831_, port_0cc0d92d_, port_4b42ea04_, port_6cf2bc2c_, port_360d45ff_, port_213bddc2_, port_0bf3d477_, port_24919790_, port_0cea4e99_, port_2374bcc1_, port_1ff44368_, port_1eaf7a9b_, port_40b0ff93_, port_67286d84_, port_4dcef735_, port_5e08959f_, port_404885f8_, port_6438f003_, RESULT, RESULT_u320, RESULT_u321, RESULT_u322, RESULT_u323, RESULT_u324, RESULT_u325, RESULT_u326, RESULT_u327, RESULT_u328, RESULT_u329, RESULT_u330, RESULT_u331, RESULT_u332, RESULT_u333, RESULT_u334, RESULT_u335, RESULT_u336, RESULT_u337, RESULT_u338, RESULT_u339, RESULT_u340, RESULT_u341, RESULT_u342, RESULT_u343, DONE);
input		CLK;
input		RESET;
input		GO;
input	[2:0]	port_42620ba7_;
input	[15:0]	port_41492b7c_;
input	[15:0]	port_34f62b85_;
input	[15:0]	port_6d2bfa2d_;
input	[31:0]	port_2e0d86cd_;
input		port_70e1f405_;
input		port_6d3af1f9_;
input		port_459c8efa_;
input		port_24157214_;
input		port_6e290ca0_;
input		port_28187583_;
input		port_5cc4abf1_;
input		port_010adde4_;
input		port_756b4eaa_;
input		port_6004d831_;
input		port_0cc0d92d_;
input		port_4b42ea04_;
input		port_6cf2bc2c_;
input		port_360d45ff_;
input		port_213bddc2_;
input		port_0bf3d477_;
input		port_24919790_;
input		port_0cea4e99_;
input		port_2374bcc1_;
input		port_1ff44368_;
input		port_1eaf7a9b_;
input		port_40b0ff93_;
input		port_67286d84_;
input		port_4dcef735_;
input		port_5e08959f_;
input		port_404885f8_;
input		port_6438f003_;
output		RESULT;
output	[2:0]	RESULT_u320;
output		RESULT_u321;
output		RESULT_u322;
output		RESULT_u323;
output		RESULT_u324;
output		RESULT_u325;
output		RESULT_u326;
output		RESULT_u327;
output		RESULT_u328;
output		RESULT_u329;
output		RESULT_u330;
output		RESULT_u331;
output		RESULT_u332;
output		RESULT_u333;
output		RESULT_u334;
output		RESULT_u335;
output		RESULT_u336;
output		RESULT_u337;
output		RESULT_u338;
output		RESULT_u339;
output		RESULT_u340;
output		RESULT_u341;
output		RESULT_u342;
output		RESULT_u343;
output		DONE;
wire		and_u391_u0;
wire signed	[15:0]	lessThan_b_signed;
wire signed	[15:0]	lessThan_a_signed;
wire		lessThan;
wire		equals;
wire signed	[15:0]	equals_b_signed;
wire signed	[15:0]	equals_a_signed;
wire		lessThan_u0;
wire	[15:0]	lessThan_u0_b_unsigned;
wire	[15:0]	lessThan_u0_a_unsigned;
wire		equals_u6;
wire	[15:0]	equals_u6_a_unsigned;
wire	[15:0]	equals_u6_b_unsigned;
wire	[15:0]	equals_u7_b_unsigned;
wire		equals_u7;
wire	[15:0]	equals_u7_a_unsigned;
wire		lessThan_u1;
wire signed	[15:0]	lessThan_u1_b_signed;
wire signed	[15:0]	lessThan_u1_a_signed;
wire		andOp;
wire	[31:0]	lessThan_u2_a_unsigned;
wire	[31:0]	lessThan_u2_b_unsigned;
wire		lessThan_u2;
wire		andOp_u0;
wire		andOp_u1;
wire	[15:0]	equals_u8_a_unsigned;
wire		equals_u8;
wire	[15:0]	equals_u8_b_unsigned;
wire		lessThan_u3;
wire signed	[15:0]	lessThan_u3_b_signed;
wire signed	[15:0]	lessThan_u3_a_signed;
wire		andOp_u2;
wire	[31:0]	lessThan_u4_a_unsigned;
wire	[31:0]	lessThan_u4_b_unsigned;
wire		lessThan_u4;
wire		andOp_u3;
wire		not_u54;
wire		andOp_u4;
wire		equals_u9;
wire	[15:0]	equals_u9_a_unsigned;
wire	[15:0]	equals_u9_b_unsigned;
wire		lessThan_u5;
wire signed	[15:0]	lessThan_u5_b_signed;
wire signed	[15:0]	lessThan_u5_a_signed;
wire		andOp_u5;
wire	[31:0]	equals_u10_a_unsigned;
wire	[31:0]	equals_u10_b_unsigned;
wire		equals_u10;
wire		andOp_u6;
wire		andOp_u7;
wire	[15:0]	equals_u11_a_unsigned;
wire		equals_u11;
wire	[15:0]	equals_u11_b_unsigned;
wire		lessThan_u6;
wire signed	[15:0]	lessThan_u6_b_signed;
wire signed	[15:0]	lessThan_u6_a_signed;
wire		andOp_u8;
wire	[31:0]	equals_u12_a_unsigned;
wire	[31:0]	equals_u12_b_unsigned;
wire		equals_u12;
wire		andOp_u9;
wire		not_u55;
wire		andOp_u10;
wire		lessThan_u7;
wire	[15:0]	lessThan_u7_b_unsigned;
wire	[15:0]	lessThan_u7_a_unsigned;
wire		lessThan_u8;
wire signed	[15:0]	lessThan_u8_b_signed;
wire signed	[15:0]	lessThan_u8_a_signed;
wire		andOp_u11;
wire		lessThan_u9;
wire	[31:0]	lessThan_u9_b_unsigned;
wire	[31:0]	lessThan_u9_a_unsigned;
wire		andOp_u12;
wire		andOp_u13;
wire		lessThan_u10;
wire	[15:0]	lessThan_u10_a_unsigned;
wire	[15:0]	lessThan_u10_b_unsigned;
wire		lessThan_u11;
wire signed	[15:0]	lessThan_u11_b_signed;
wire signed	[15:0]	lessThan_u11_a_signed;
wire		andOp_u14;
wire	[31:0]	lessThan_u12_a_unsigned;
wire		lessThan_u12;
wire	[31:0]	lessThan_u12_b_unsigned;
wire		andOp_u15;
wire		not_u56;
wire		andOp_u16;
wire	[15:0]	lessThan_u13_a_unsigned;
wire	[15:0]	lessThan_u13_b_unsigned;
wire		lessThan_u13;
wire	[31:0]	equals_u13_a_unsigned;
wire		equals_u13;
wire	[31:0]	equals_u13_b_unsigned;
wire		andOp_u17;
wire		andOp_u18;
wire		lessThan_u14;
wire	[15:0]	lessThan_u14_a_unsigned;
wire	[15:0]	lessThan_u14_b_unsigned;
wire		equals_u14;
wire	[31:0]	equals_u14_b_unsigned;
wire	[31:0]	equals_u14_a_unsigned;
wire		andOp_u19;
wire		not_u57;
wire		andOp_u20;
wire		equals_u15;
wire	[15:0]	equals_u15_b_unsigned;
wire	[15:0]	equals_u15_a_unsigned;
wire	[31:0]	lessThan_u15_a_unsigned;
wire	[31:0]	lessThan_u15_b_unsigned;
wire		lessThan_u15;
wire		andOp_u21;
wire		andOp_u22;
wire	[15:0]	equals_u16_b_unsigned;
wire	[15:0]	equals_u16_a_unsigned;
wire		equals_u16;
wire	[31:0]	lessThan_u16_a_unsigned;
wire	[31:0]	lessThan_u16_b_unsigned;
wire		lessThan_u16;
wire		andOp_u23;
wire		not_u58;
wire		andOp_u24;
wire		equals_u17;
wire	[15:0]	equals_u17_b_unsigned;
wire	[15:0]	equals_u17_a_unsigned;
wire	[31:0]	equals_u18_b_unsigned;
wire	[31:0]	equals_u18_a_unsigned;
wire		equals_u18;
wire		andOp_u25;
wire		andOp_u26;
wire	[15:0]	equals_u19_b_unsigned;
wire	[15:0]	equals_u19_a_unsigned;
wire		equals_u19;
wire	[31:0]	equals_u20_b_unsigned;
wire		equals_u20;
wire	[31:0]	equals_u20_a_unsigned;
wire		andOp_u27;
wire		not_u59;
wire		andOp_u28;
wire	[15:0]	equals_u21_b_unsigned;
wire	[15:0]	equals_u21_a_unsigned;
wire		equals_u21;
wire signed	[15:0]	equals_u22_a_signed;
wire		equals_u22;
wire signed	[15:0]	equals_u22_b_signed;
wire		andOp_u29;
wire	[31:0]	equals_u23_b_unsigned;
wire		equals_u23;
wire	[31:0]	equals_u23_a_unsigned;
wire		andOp_u30;
wire		andOp_u31;
wire	[15:0]	equals_u24_b_unsigned;
wire		equals_u24;
wire	[15:0]	equals_u24_a_unsigned;
wire signed	[15:0]	equals_u25_b_signed;
wire signed	[15:0]	equals_u25_a_signed;
wire		equals_u25;
wire		andOp_u32;
wire	[31:0]	equals_u26_a_unsigned;
wire	[31:0]	equals_u26_b_unsigned;
wire		equals_u26;
wire		andOp_u33;
wire		not_u60;
wire		andOp_u34;
wire	[15:0]	lessThan_u17_a_unsigned;
wire	[15:0]	lessThan_u17_b_unsigned;
wire		lessThan_u17;
wire		equals_u27;
wire	[31:0]	equals_u27_a_unsigned;
wire	[31:0]	equals_u27_b_unsigned;
wire		andOp_u35;
wire		andOp_u36;
wire		lessThan_u18;
wire	[15:0]	lessThan_u18_a_unsigned;
wire	[15:0]	lessThan_u18_b_unsigned;
wire		equals_u28;
wire	[31:0]	equals_u28_a_unsigned;
wire	[31:0]	equals_u28_b_unsigned;
wire		andOp_u37;
wire		not_u61;
wire		andOp_u38;
wire	[15:0]	equals_u29_b_unsigned;
wire	[15:0]	equals_u29_a_unsigned;
wire		equals_u29;
wire	[31:0]	equals_u30_a_unsigned;
wire	[31:0]	equals_u30_b_unsigned;
wire		equals_u30;
wire		andOp_u39;
wire		andOp_u40;
wire	[15:0]	equals_u31_a_unsigned;
wire		equals_u31;
wire	[15:0]	equals_u31_b_unsigned;
wire	[31:0]	equals_u32_a_unsigned;
wire		equals_u32;
wire	[31:0]	equals_u32_b_unsigned;
wire		andOp_u41;
wire		not_u62;
wire		andOp_u42;
wire signed	[31:0]	equals_u33_b_signed;
wire signed	[31:0]	equals_u33_a_signed;
wire		equals_u33;
wire		and_u392_u0;
wire		not_u63_u0;
wire		and_u393_u0;
wire		andOp_u43;
wire		not_u64_u0;
wire		and_u394_u0;
wire		and_u395_u0;
wire		simplePinWrite;
wire		and_u396_u0;
wire		not_u65_u0;
wire		and_u397_u0;
wire		simplePinWrite_u74;
wire		and_u398_u0;
wire		and_u399_u0;
wire		or_u86_u0;
wire	[2:0]	mux_u28;
wire		and_u400_u0;
wire		and_u401_u0;
wire signed	[31:0]	equals_u34_a_signed;
wire signed	[31:0]	equals_u34_b_signed;
wire		equals_u34;
wire		and_u402_u0;
wire		not_u66_u0;
wire		and_u403_u0;
wire		and_u404_u0;
wire		not_u67_u0;
wire		and_u405_u0;
wire		and_u406_u0;
wire		and_u407_u0;
wire		not_u68_u0;
wire		simplePinWrite_u75;
reg		reg_3a1f45fa_u0=1'h0;
reg		reg_75145b92_u0=1'h0;
reg		reg_747e49b6_u0=1'h0;
wire		and_u408_u0;
reg		reg_33c17034_u0=1'h0;
wire		and_u409_u0;
reg		reg_33c17034_result_delayed_u0=1'h0;
reg		reg_3a1f45fa_result_delayed_u0=1'h0;
reg		reg_75145b92_result_delayed_u0=1'h0;
wire		or_u87_u0;
reg		reg_66d1b020_u0=1'h0;
wire		and_u410_u0;
wire		or_u88_u0;
wire		and_u411_u0;
reg		reg_1b67eb07_u0=1'h0;
wire		and_u412_u0;
wire		and_u413_u0;
wire		or_u89_u0;
wire signed	[31:0]	equals_u35_a_signed;
wire signed	[31:0]	equals_u35_b_signed;
wire		equals_u35;
wire		and_u414_u0;
wire		not_u69_u0;
wire		and_u415_u0;
wire		andOp_u44;
wire		not_u70_u0;
wire		and_u416_u0;
wire		and_u417_u0;
wire		and_u418_u0;
wire		not_u71_u0;
wire		and_u419_u0;
wire		simplePinWrite_u76;
wire		and_u420_u0;
reg		reg_179dcff8_u0=1'h0;
reg		reg_7d7c20fb_u0=1'h0;
wire		and_u421_u0;
reg		reg_0322b1ca_u0=1'h0;
reg		reg_38422e0b_u0=1'h0;
wire		or_u90_u0;
reg		and_delayed_u4=1'h0;
reg		reg_7d7c20fb_result_delayed_u0=1'h0;
reg		reg_179dcff8_result_delayed_u0=1'h0;
wire		andOp_u45;
wire		and_u422_u0;
wire		not_u72_u0;
wire		and_u423_u0;
wire		and_u424_u0;
wire		and_u425_u0;
wire		not_u73_u0;
wire		simplePinWrite_u77;
reg		reg_6f660aa7_u0=1'h0;
reg		reg_1a2c6ea5_u0=1'h0;
wire		or_u91_u0;
wire		and_u426_u0;
reg		reg_6f660aa7_result_delayed_u0=1'h0;
reg		reg_2e392276_u0=1'h0;
reg		reg_115cba2e_u0=1'h0;
wire		and_u427_u0;
reg		reg_1a2c6ea5_result_delayed_u0=1'h0;
reg		reg_6f660aa7_result_delayed_result_delayed_u0=1'h0;
wire		and_u428_u0;
wire		and_u429_u0;
reg		and_delayed_u5_u0=1'h0;
wire		or_u92_u0;
wire		or_u93_u0;
wire	[2:0]	mux_u29_u0;
wire		and_u430_u0;
wire		or_u94_u0;
wire		and_u431_u0;
reg		reg_3f285a69_u0=1'h0;
wire		and_u432_u0;
wire		and_u433_u0;
wire		or_u95_u0;
wire signed	[31:0]	equals_u36_a_signed;
wire		equals_u36;
wire signed	[31:0]	equals_u36_b_signed;
wire		not_u74_u0;
wire		and_u434_u0;
wire		and_u435_u0;
wire		andOp_u46;
wire		and_u436_u0;
wire		and_u437_u0;
wire		not_u75_u0;
wire		and_u438_u0;
wire		not_u76_u0;
wire		and_u439_u0;
wire		simplePinWrite_u78;
wire		or_u96_u0;
reg		reg_4fb73053_u0=1'h0;
wire		and_u440_u0;
reg		reg_6a7d31d4_u0=1'h0;
reg		and_delayed_u6_u0=1'h0;
reg		reg_63ede03c_u0=1'h0;
wire		and_u441_u0;
reg		reg_4fb73053_result_delayed_u0=1'h0;
reg		reg_6a7d31d4_result_delayed_u0=1'h0;
reg		reg_6a7d31d4_result_delayed_result_delayed_u0=1'h0;
wire		andOp_u47;
wire		not_u77_u0;
wire		and_u442_u0;
wire		and_u443_u0;
wire		and_u444_u0;
wire		not_u78_u0;
wire		and_u445_u0;
wire		simplePinWrite_u79;
wire		and_u446_u0;
reg		reg_4dff0c7d_u0=1'h0;
reg		reg_4dff0c7d_result_delayed_u0=1'h0;
wire		and_u447_u0;
wire		or_u97_u0;
reg		reg_4056b2dd_u0=1'h0;
reg		reg_0da41b16_u0=1'h0;
reg		reg_4dff0c7d_result_delayed_result_delayed_u0=1'h0;
reg		and_delayed_u7_u0=1'h0;
reg		reg_4056b2dd_result_delayed_u0=1'h0;
wire		not_u79_u0;
wire		and_u448_u0;
wire		and_u449_u0;
wire		not_u80_u0;
wire		and_u450_u0;
wire		and_u451_u0;
wire		simplePinWrite_u80;
reg		reg_39b080d6_u0=1'h0;
reg		reg_54f4b899_u0=1'h0;
reg		reg_54f4b899_result_delayed_u0=1'h0;
reg		reg_66a4207d_u0=1'h0;
wire		and_u452_u0;
reg		reg_7c85adb8_u0=1'h0;
wire		or_u98_u0;
reg		reg_54f4b899_result_delayed_result_delayed_u0=1'h0;
wire		and_u453_u0;
wire		and_u454_u0;
wire		and_u455_u0;
wire		not_u81_u0;
wire		and_u456_u0;
wire		and_u457_u0;
wire		not_u82_u0;
wire		simplePinWrite_u81;
wire		and_u458_u0;
reg		reg_67690009_u0=1'h0;
reg		reg_2eb38cd6_u0=1'h0;
wire		or_u99_u0;
reg		and_delayed_u8_u0=1'h0;
wire		and_u459_u0;
reg		reg_2eb38cd6_result_delayed_u0=1'h0;
reg		reg_67690009_result_delayed_u0=1'h0;
reg		and_delayed_u9_u0=1'h0;
wire		and_u460_u0;
reg		and_delayed_u10_u0=1'h0;
wire		or_u100_u0;
wire		and_u461_u0;
wire		or_u101_u0;
wire		and_u462_u0;
wire		and_u463_u0;
wire		or_u102_u0;
wire		and_u464_u0;
wire		or_u103_u0;
wire		or_u104_u0;
wire		and_u465_u0;
wire		or_u105_u0;
wire		and_u466_u0;
wire		and_u467_u0;
wire		or_u106_u0;
reg		reg_4e472843_u0=1'h0;
wire		and_u468_u0;
wire		and_u469_u0;
wire		or_u107_u0;
wire signed	[31:0]	equals_u37_a_signed;
wire signed	[31:0]	equals_u37_b_signed;
wire		equals_u37;
wire		and_u470_u0;
wire		and_u471_u0;
wire		not_u83_u0;
wire		andOp_u48;
wire		and_u472_u0;
wire		not_u84_u0;
wire		and_u473_u0;
wire		not_u85_u0;
wire		and_u474_u0;
wire		and_u475_u0;
wire		simplePinWrite_u82;
reg		reg_6e3a0db9_u0=1'h0;
reg		reg_43d57d30_u0=1'h0;
reg		reg_4d5434d2_u0=1'h0;
reg		reg_5bff6a34_u0=1'h0;
reg		reg_5bff6a34_result_delayed_u0=1'h0;
wire		or_u108_u0;
wire		and_u476_u0;
wire		and_u477_u0;
reg		reg_5bff6a34_result_delayed_result_delayed_u0=1'h0;
reg		reg_4d5434d2_result_delayed_u0=1'h0;
wire		andOp_u49;
wire		and_u478_u0;
wire		not_u86_u0;
wire		and_u479_u0;
wire		not_u87_u0;
wire		and_u480_u0;
wire		and_u481_u0;
wire		simplePinWrite_u83;
wire		or_u109_u0;
reg		reg_7b478222_u0=1'h0;
reg		reg_2e3fd957_u0=1'h0;
reg		reg_48ed0ea7_u0=1'h0;
wire		and_u482_u0;
reg		reg_48ed0ea7_result_delayed_u0=1'h0;
reg		reg_6b6f3e79_u0=1'h0;
reg		reg_2e3fd957_result_delayed_u0=1'h0;
wire		and_u483_u0;
reg		reg_2e3fd957_result_delayed_result_delayed_u0=1'h0;
wire		not_u88_u0;
wire		and_u484_u0;
wire		and_u485_u0;
wire		not_u89_u0;
wire		and_u486_u0;
wire		and_u487_u0;
wire		simplePinWrite_u84;
reg		reg_6d9aed1d_u0=1'h0;
reg		reg_5afb3453_u0=1'h0;
wire		and_u488_u0;
reg		reg_1c6adbe7_u0=1'h0;
reg		reg_6d9aed1d_result_delayed_u0=1'h0;
reg		reg_1decc03f_u0=1'h0;
reg		reg_1decc03f_result_delayed_u0=1'h0;
wire		and_u489_u0;
wire		or_u110_u0;
wire		not_u90_u0;
wire		and_u490_u0;
wire		and_u491_u0;
wire		and_u492_u0;
wire		not_u91_u0;
wire		and_u493_u0;
wire		simplePinWrite_u85;
reg		reg_2b6f460f_u0=1'h0;
wire		and_u494_u0;
wire		and_u495_u0;
reg		reg_2b6f460f_result_delayed_u0=1'h0;
wire		or_u111_u0;
reg		reg_2b6f460f_result_delayed_result_delayed_u0=1'h0;
reg		reg_4138b0a0_u0=1'h0;
reg		and_delayed_u11_u0=1'h0;
reg		and_delayed_u12_u0=1'h0;
wire		andOp_u50;
wire		and_u496_u0;
wire		not_u92_u0;
wire		and_u497_u0;
wire		and_u498_u0;
wire		and_u499_u0;
wire		not_u93_u0;
wire		simplePinWrite_u86;
reg		reg_5475b2b5_u0=1'h0;
wire		and_u500_u0;
wire		and_u501_u0;
reg		reg_7c3d02d5_u0=1'h0;
reg		reg_7c3d02d5_result_delayed_u0=1'h0;
reg		reg_424c04bc_u0=1'h0;
reg		reg_424c04bc_result_delayed_u0=1'h0;
reg		reg_7c3d02d5_result_delayed_result_delayed_u0=1'h0;
reg		and_delayed_u13_u0=1'h0;
wire		or_u112_u0;
wire		andOp_u51;
wire		not_u94_u0;
wire		and_u502_u0;
wire		and_u503_u0;
wire		and_u504_u0;
wire		not_u95_u0;
wire		and_u505_u0;
wire		simplePinWrite_u87;
reg		reg_71b65551_u0=1'h0;
reg		reg_5557b19e_u0=1'h0;
reg		reg_117d0bd6_u0=1'h0;
wire		or_u113_u0;
wire		and_u506_u0;
wire		and_u507_u0;
reg		and_delayed_u14_u0=1'h0;
reg		and_delayed_result_delayed_u0=1'h0;
reg		reg_71b65551_result_delayed_u0=1'h0;
reg		and_delayed_result_delayed_result_delayed_u0=1'h0;
wire		and_u508_u0;
wire		and_u509_u0;
wire		not_u96_u0;
wire		and_u510_u0;
wire		not_u97_u0;
wire		and_u511_u0;
wire		simplePinWrite_u88;
reg		reg_04f3c4f4_u0=1'h0;
reg		reg_76e06d48_u0=1'h0;
reg		reg_7d698f03_u0=1'h0;
wire		and_u512_u0;
reg		reg_7d698f03_result_delayed_u0=1'h0;
reg		and_delayed_u15_u0=1'h0;
reg		reg_04f3c4f4_result_delayed_u0=1'h0;
wire		or_u114_u0;
wire		and_u513_u0;
wire		and_u514_u0;
wire		not_u98_u0;
wire		and_u515_u0;
wire		and_u516_u0;
wire		and_u517_u0;
wire		not_u99_u0;
wire		simplePinWrite_u89;
reg		reg_5b4fb5ce_u0=1'h0;
wire		and_u518_u0;
reg		reg_52c1fee5_u0=1'h0;
reg		reg_1ccb0e6e_u0=1'h0;
reg		and_delayed_u16_u0=1'h0;
wire		or_u115_u0;
reg		reg_26f8fd95_u0=1'h0;
wire		and_u519_u0;
reg		reg_5b4fb5ce_result_delayed_u0=1'h0;
wire		and_u520_u0;
wire		or_u116_u0;
reg		and_delayed_u17_u0=1'h0;
wire		and_u521_u0;
wire		and_u522_u0;
wire		and_u523_u0;
wire		or_u117_u0;
wire		or_u118_u0;
wire		or_u119_u0;
wire		or_u120_u0;
wire		and_u524_u0;
wire		and_u525_u0;
wire		and_u526_u0;
wire		or_u121_u0;
wire		or_u122_u0;
wire		and_u527_u0;
wire	[2:0]	mux_u30_u0;
wire		or_u123_u0;
wire		and_u528_u0;
wire		or_u124_u0;
wire		and_u529_u0;
wire		and_u530_u0;
wire		and_u531_u0;
wire		or_u125_u0;
wire	[2:0]	mux_u31_u0;
wire		or_u126_u0;
wire		and_u532_u0;
wire		and_u533_u0;
wire		or_u127_u0;
wire		or_u128_u0;
wire	[2:0]	mux_u32_u0;
wire		and_u534_u0;
wire		and_u535_u0;
wire		or_u129_u0;
wire	[2:0]	mux_u33_u0;
wire		or_u130_u0;
wire		or_u131_u0;
wire		and_u536_u0;
wire		and_u537_u0;
reg		and_delayed_u18_u0=1'h0;
wire signed	[31:0]	equals_u38_a_signed;
wire signed	[31:0]	equals_u38_b_signed;
wire		equals_u38;
wire		not_u100_u0;
wire		and_u538_u0;
wire		and_u539_u0;
wire		andOp_u52;
wire		and_u540_u0;
wire		not_u101_u0;
wire		and_u541_u0;
wire		not_u102_u0;
wire		and_u542_u0;
wire		and_u543_u0;
wire		simplePinWrite_u90;
reg		reg_60e797c7_u0=1'h0;
wire		or_u132_u0;
reg		reg_14bc455b_u0=1'h0;
reg		reg_14bc455b_result_delayed_u0=1'h0;
wire		and_u544_u0;
reg		and_delayed_u19_u0=1'h0;
wire		and_u545_u0;
reg		and_delayed_u20_u0=1'h0;
reg		reg_01c7fa9c_u0=1'h0;
reg		and_delayed_result_delayed_u1_u0=1'h0;
wire		andOp_u53;
wire		and_u546_u0;
wire		and_u547_u0;
wire		not_u103_u0;
wire		and_u548_u0;
wire		and_u549_u0;
wire		not_u104_u0;
wire		simplePinWrite_u91;
wire		and_u550_u0;
reg		reg_7b1e075a_u0=1'h0;
reg		reg_37e60342_u0=1'h0;
reg		reg_0834cf70_u0=1'h0;
reg		reg_37e60342_result_delayed_u0=1'h0;
reg		reg_7b1e075a_result_delayed_u0=1'h0;
wire		and_u551_u0;
reg		reg_7b1e075a_result_delayed_result_delayed_u0=1'h0;
wire		or_u133_u0;
reg		and_delayed_u21_u0=1'h0;
wire		and_u552_u0;
wire		and_u553_u0;
wire		not_u105_u0;
wire		and_u554_u0;
wire		and_u555_u0;
wire		not_u106_u0;
wire		simplePinWrite_u92;
reg		reg_2b889e88_u0=1'h0;
reg		reg_3fd6f110_u0=1'h0;
wire		and_u556_u0;
reg		reg_33af66c3_u0=1'h0;
reg		reg_2b889e88_result_delayed_u0=1'h0;
wire		and_u557_u0;
reg		and_delayed_u22_u0=1'h0;
wire		or_u134_u0;
reg		reg_3fd6f110_result_delayed_u0=1'h0;
wire		not_u107_u0;
wire		and_u558_u0;
wire		and_u559_u0;
wire		and_u560_u0;
wire		and_u561_u0;
wire		not_u108_u0;
wire		simplePinWrite_u93;
reg		reg_49ed7469_u0=1'h0;
reg		reg_575d09b8_u0=1'h0;
wire		and_u562_u0;
wire		and_u563_u0;
reg		reg_6efc1130_u0=1'h0;
reg		reg_49ed7469_result_delayed_u0=1'h0;
wire		or_u135_u0;
reg		reg_49ed7469_result_delayed_result_delayed_u0=1'h0;
reg		and_delayed_u23_u0=1'h0;
wire		and_u564_u0;
wire		not_u109_u0;
wire		and_u565_u0;
wire		and_u566_u0;
wire		and_u567_u0;
wire		not_u110_u0;
wire		simplePinWrite_u94;
wire		and_u568_u0;
wire		and_u569_u0;
reg		and_delayed_u24_u0=1'h0;
reg		reg_1723f867_u0=1'h0;
reg		reg_11292ccc_u0=1'h0;
reg		reg_11292ccc_result_delayed_u0=1'h0;
reg		and_delayed_u25_u0=1'h0;
wire		or_u136_u0;
reg		reg_11292ccc_result_delayed_result_delayed_u0=1'h0;
wire		and_u570_u0;
wire		and_u571_u0;
wire		not_u111_u0;
wire		not_u112_u0;
wire		and_u572_u0;
wire		and_u573_u0;
wire		simplePinWrite_u95;
reg		reg_64e07a44_u0=1'h0;
reg		reg_23dba81c_u0=1'h0;
reg		reg_23dba81c_result_delayed_u0=1'h0;
reg		reg_15bcd7f0_u0=1'h0;
wire		and_u574_u0;
reg		reg_53451f0b_u0=1'h0;
wire		and_u575_u0;
reg		reg_23dba81c_result_delayed_result_delayed_u0=1'h0;
wire		or_u137_u0;
reg		reg_106be70b_u0=1'h0;
wire		and_u576_u0;
wire		or_u138_u0;
wire		and_u577_u0;
wire		or_u139_u0;
wire		and_u578_u0;
wire		and_u579_u0;
wire		or_u140_u0;
wire		and_u580_u0;
wire		and_u581_u0;
wire		or_u141_u0;
wire	[2:0]	mux_u34_u0;
wire		or_u142_u0;
wire		and_u582_u0;
wire		and_u583_u0;
wire	[2:0]	mux_u35_u0;
wire		or_u143_u0;
wire		or_u144_u0;
wire		and_u584_u0;
wire		and_u585_u0;
wire	[2:0]	mux_u36_u0;
wire		or_u145_u0;
wire		or_u146_u0;
wire		and_u586_u0;
wire		or_u147_u0;
wire	[2:0]	mux_u37_u0;
wire		and_u587_u0;
wire		or_u148_u0;
wire		or_u149_u0;
wire		and_u588_u0;
reg		reg_1032f60e_u0=1'h0;
wire		and_u589_u0;
wire signed	[31:0]	equals_u39_a_signed;
wire signed	[31:0]	equals_u39_b_signed;
wire		equals_u39;
wire		and_u590_u0;
wire		and_u591_u0;
wire		not_u113_u0;
wire		and_u592_u0;
wire		not_u114_u0;
wire		and_u593_u0;
wire		and_u594_u0;
wire		and_u595_u0;
wire		not_u115_u0;
wire		simplePinWrite_u96;
reg		reg_631bc458_u0=1'h0;
reg		reg_67355df6_u0=1'h0;
wire		or_u150_u0;
reg		reg_07f5313f_u0=1'h0;
reg		reg_789509d9_u0=1'h0;
wire		and_u596_u0;
reg		reg_631bc458_result_delayed_u0=1'h0;
wire		and_u597_u0;
reg		reg_789509d9_result_delayed_u0=1'h0;
wire		not_u116_u0;
wire		and_u598_u0;
wire		and_u599_u0;
wire		and_u600_u0;
wire		and_u601_u0;
wire		not_u117_u0;
wire		simplePinWrite_u97;
reg		reg_45853e06_u0=1'h0;
reg		reg_45853e06_result_delayed_u0=1'h0;
wire		and_u602_u0;
reg		reg_00fcf046_u0=1'h0;
wire		or_u151_u0;
wire		and_u603_u0;
reg		and_delayed_u26_u0=1'h0;
reg		and_delayed_u27_u0=1'h0;
reg		reg_45853e06_result_delayed_result_delayed_u0=1'h0;
wire		and_u604_u0;
wire		not_u118_u0;
wire		and_u605_u0;
wire		and_u606_u0;
wire		not_u119_u0;
wire		and_u607_u0;
wire		simplePinWrite_u98;
reg		reg_4b138e52_u0=1'h0;
reg		reg_6bcd16e4_u0=1'h0;
wire		and_u608_u0;
reg		reg_36c01350_u0=1'h0;
reg		reg_36c01350_result_delayed_u0=1'h0;
reg		and_delayed_u28_u0=1'h0;
wire		and_u609_u0;
wire		or_u152_u0;
reg		reg_4b138e52_result_delayed_u0=1'h0;
wire		and_u610_u0;
wire		not_u120_u0;
wire		and_u611_u0;
wire		and_u612_u0;
wire		and_u613_u0;
wire		not_u121_u0;
wire		simplePinWrite_u99;
wire		and_u614_u0;
reg		and_delayed_u29_u0=1'h0;
reg		and_delayed_result_delayed_u2_u0=1'h0;
reg		reg_265a004b_u0=1'h0;
reg		reg_265a004b_result_delayed_u0=1'h0;
reg		reg_60ff05ab_u0=1'h0;
wire		and_u615_u0;
reg		and_delayed_result_delayed_result_delayed_u1_u0=1'h0;
wire		or_u153_u0;
wire		and_u616_u0;
reg		reg_20083bde_u0=1'h0;
wire		and_u617_u0;
wire		or_u154_u0;
wire		and_u618_u0;
wire		or_u155_u0;
wire		and_u619_u0;
wire		or_u156_u0;
wire		and_u620_u0;
wire		or_u157_u0;
wire		and_u621_u0;
wire		or_u158_u0;
wire	[2:0]	mux_u38_u0;
wire		or_u159_u0;
wire		and_u622_u0;
wire		or_u160_u0;
wire	[2:0]	mux_u39_u0;
wire		and_u623_u0;
wire		and_u624_u0;
wire		and_u625_u0;
wire		or_u161_u0;
reg		and_delayed_u30_u0=1'h0;
wire		midLeft2_go_merge;
wire		midLeft1_go_merge;
wire		midLeftNoConsume2_go_merge;
wire		midLeftNoConsume1_go_merge;
wire		scoreboard_45f1cb9d_and;
reg		scoreboard_45f1cb9d_reg0=1'h0;
wire		scoreboard_45f1cb9d_resOr3;
wire		bus_384ef3c0_;
wire		scoreboard_45f1cb9d_resOr4;
wire		scoreboard_45f1cb9d_resOr0;
reg		scoreboard_45f1cb9d_reg1=1'h0;
reg		scoreboard_45f1cb9d_reg5=1'h0;
reg		scoreboard_45f1cb9d_reg3=1'h0;
wire		scoreboard_45f1cb9d_resOr2;
reg		scoreboard_45f1cb9d_reg4=1'h0;
wire		scoreboard_45f1cb9d_resOr1;
reg		scoreboard_45f1cb9d_reg2=1'h0;
wire		scoreboard_45f1cb9d_resOr5;
wire	[2:0]	mux_u40_u0;
wire		or_u162_u0;
wire		or_u163_u0;
reg		reg_45547147_u0=1'h0;
wire	[2:0]	mux_u41_u0;
wire		or_u164_u0;
reg		reg_45547147_result_delayed_u0=1'h0;
assign and_u391_u0=or_u163_u0&or_u163_u0;
assign lessThan_a_signed=port_41492b7c_;
assign lessThan_b_signed=16'h103;
assign lessThan=lessThan_a_signed<lessThan_b_signed;
assign equals_a_signed=port_41492b7c_;
assign equals_b_signed=16'h103;
assign equals=equals_a_signed==equals_b_signed;
assign lessThan_u0_a_unsigned=port_34f62b85_;
assign lessThan_u0_b_unsigned=16'hff;
assign lessThan_u0=lessThan_u0_a_unsigned<lessThan_u0_b_unsigned;
assign equals_u6_a_unsigned=port_34f62b85_;
assign equals_u6_b_unsigned=16'hff;
assign equals_u6=equals_u6_a_unsigned==equals_u6_b_unsigned;
assign equals_u7_a_unsigned=port_34f62b85_;
assign equals_u7_b_unsigned=16'h0;
assign equals_u7=equals_u7_a_unsigned==equals_u7_b_unsigned;
assign lessThan_u1_a_signed=port_6d2bfa2d_;
assign lessThan_u1_b_signed=16'h1ff;
assign lessThan_u1=lessThan_u1_a_signed<lessThan_u1_b_signed;
assign andOp=equals_u7&lessThan_u1;
assign lessThan_u2_a_unsigned=port_2e0d86cd_;
assign lessThan_u2_b_unsigned=32'h20000;
assign lessThan_u2=lessThan_u2_a_unsigned<lessThan_u2_b_unsigned;
assign andOp_u0=andOp&lessThan_u2;
assign andOp_u1=andOp_u0&port_70e1f405_;
assign equals_u8_a_unsigned=port_34f62b85_;
assign equals_u8_b_unsigned=16'h0;
assign equals_u8=equals_u8_a_unsigned==equals_u8_b_unsigned;
assign lessThan_u3_a_signed=port_6d2bfa2d_;
assign lessThan_u3_b_signed=16'h1ff;
assign lessThan_u3=lessThan_u3_a_signed<lessThan_u3_b_signed;
assign andOp_u2=equals_u8&lessThan_u3;
assign lessThan_u4_a_unsigned=port_2e0d86cd_;
assign lessThan_u4_b_unsigned=32'h20000;
assign lessThan_u4=lessThan_u4_a_unsigned<lessThan_u4_b_unsigned;
assign andOp_u3=andOp_u2&lessThan_u4;
assign not_u54=!port_70e1f405_;
assign andOp_u4=andOp_u3&not_u54;
assign equals_u9_a_unsigned=port_34f62b85_;
assign equals_u9_b_unsigned=16'h0;
assign equals_u9=equals_u9_a_unsigned==equals_u9_b_unsigned;
assign lessThan_u5_a_signed=port_6d2bfa2d_;
assign lessThan_u5_b_signed=16'h1ff;
assign lessThan_u5=lessThan_u5_a_signed<lessThan_u5_b_signed;
assign andOp_u5=equals_u9&lessThan_u5;
assign equals_u10_a_unsigned=port_2e0d86cd_;
assign equals_u10_b_unsigned=32'h20000;
assign equals_u10=equals_u10_a_unsigned==equals_u10_b_unsigned;
assign andOp_u6=andOp_u5&equals_u10;
assign andOp_u7=andOp_u6&port_70e1f405_;
assign equals_u11_a_unsigned=port_34f62b85_;
assign equals_u11_b_unsigned=16'h0;
assign equals_u11=equals_u11_a_unsigned==equals_u11_b_unsigned;
assign lessThan_u6_a_signed=port_6d2bfa2d_;
assign lessThan_u6_b_signed=16'h1ff;
assign lessThan_u6=lessThan_u6_a_signed<lessThan_u6_b_signed;
assign andOp_u8=equals_u11&lessThan_u6;
assign equals_u12_a_unsigned=port_2e0d86cd_;
assign equals_u12_b_unsigned=32'h20000;
assign equals_u12=equals_u12_a_unsigned==equals_u12_b_unsigned;
assign andOp_u9=andOp_u8&equals_u12;
assign not_u55=!port_70e1f405_;
assign andOp_u10=andOp_u9&not_u55;
assign lessThan_u7_a_unsigned=port_34f62b85_;
assign lessThan_u7_b_unsigned=16'hff;
assign lessThan_u7=lessThan_u7_a_unsigned<lessThan_u7_b_unsigned;
assign lessThan_u8_a_signed=port_6d2bfa2d_;
assign lessThan_u8_b_signed=16'h1ff;
assign lessThan_u8=lessThan_u8_a_signed<lessThan_u8_b_signed;
assign andOp_u11=lessThan_u7&lessThan_u8;
assign lessThan_u9_a_unsigned=port_2e0d86cd_;
assign lessThan_u9_b_unsigned=32'h20000;
assign lessThan_u9=lessThan_u9_a_unsigned<lessThan_u9_b_unsigned;
assign andOp_u12=andOp_u11&lessThan_u9;
assign andOp_u13=andOp_u12&port_70e1f405_;
assign lessThan_u10_a_unsigned=port_34f62b85_;
assign lessThan_u10_b_unsigned=16'hff;
assign lessThan_u10=lessThan_u10_a_unsigned<lessThan_u10_b_unsigned;
assign lessThan_u11_a_signed=port_6d2bfa2d_;
assign lessThan_u11_b_signed=16'h1ff;
assign lessThan_u11=lessThan_u11_a_signed<lessThan_u11_b_signed;
assign andOp_u14=lessThan_u10&lessThan_u11;
assign lessThan_u12_a_unsigned=port_2e0d86cd_;
assign lessThan_u12_b_unsigned=32'h20000;
assign lessThan_u12=lessThan_u12_a_unsigned<lessThan_u12_b_unsigned;
assign andOp_u15=andOp_u14&lessThan_u12;
assign not_u56=!port_70e1f405_;
assign andOp_u16=andOp_u15&not_u56;
assign lessThan_u13_a_unsigned=port_34f62b85_;
assign lessThan_u13_b_unsigned=16'hff;
assign lessThan_u13=lessThan_u13_a_unsigned<lessThan_u13_b_unsigned;
assign equals_u13_a_unsigned=port_2e0d86cd_;
assign equals_u13_b_unsigned=32'h20000;
assign equals_u13=equals_u13_a_unsigned==equals_u13_b_unsigned;
assign andOp_u17=lessThan_u13&equals_u13;
assign andOp_u18=andOp_u17&port_70e1f405_;
assign lessThan_u14_a_unsigned=port_34f62b85_;
assign lessThan_u14_b_unsigned=16'hff;
assign lessThan_u14=lessThan_u14_a_unsigned<lessThan_u14_b_unsigned;
assign equals_u14_a_unsigned=port_2e0d86cd_;
assign equals_u14_b_unsigned=32'h20000;
assign equals_u14=equals_u14_a_unsigned==equals_u14_b_unsigned;
assign andOp_u19=lessThan_u14&equals_u14;
assign not_u57=!port_70e1f405_;
assign andOp_u20=andOp_u19&not_u57;
assign equals_u15_a_unsigned=port_34f62b85_;
assign equals_u15_b_unsigned=16'hff;
assign equals_u15=equals_u15_a_unsigned==equals_u15_b_unsigned;
assign lessThan_u15_a_unsigned=port_2e0d86cd_;
assign lessThan_u15_b_unsigned=32'h20000;
assign lessThan_u15=lessThan_u15_a_unsigned<lessThan_u15_b_unsigned;
assign andOp_u21=equals_u15&lessThan_u15;
assign andOp_u22=andOp_u21&port_70e1f405_;
assign equals_u16_a_unsigned=port_34f62b85_;
assign equals_u16_b_unsigned=16'hff;
assign equals_u16=equals_u16_a_unsigned==equals_u16_b_unsigned;
assign lessThan_u16_a_unsigned=port_2e0d86cd_;
assign lessThan_u16_b_unsigned=32'h20000;
assign lessThan_u16=lessThan_u16_a_unsigned<lessThan_u16_b_unsigned;
assign andOp_u23=equals_u16&lessThan_u16;
assign not_u58=!port_70e1f405_;
assign andOp_u24=andOp_u23&not_u58;
assign equals_u17_a_unsigned=port_34f62b85_;
assign equals_u17_b_unsigned=16'hff;
assign equals_u17=equals_u17_a_unsigned==equals_u17_b_unsigned;
assign equals_u18_a_unsigned=port_2e0d86cd_;
assign equals_u18_b_unsigned=32'h20000;
assign equals_u18=equals_u18_a_unsigned==equals_u18_b_unsigned;
assign andOp_u25=equals_u17&equals_u18;
assign andOp_u26=andOp_u25&port_70e1f405_;
assign equals_u19_a_unsigned=port_34f62b85_;
assign equals_u19_b_unsigned=16'hff;
assign equals_u19=equals_u19_a_unsigned==equals_u19_b_unsigned;
assign equals_u20_a_unsigned=port_2e0d86cd_;
assign equals_u20_b_unsigned=32'h20000;
assign equals_u20=equals_u20_a_unsigned==equals_u20_b_unsigned;
assign andOp_u27=equals_u19&equals_u20;
assign not_u59=!port_70e1f405_;
assign andOp_u28=andOp_u27&not_u59;
assign equals_u21_a_unsigned=port_34f62b85_;
assign equals_u21_b_unsigned=16'h0;
assign equals_u21=equals_u21_a_unsigned==equals_u21_b_unsigned;
assign equals_u22_a_signed=port_6d2bfa2d_;
assign equals_u22_b_signed=16'h1ff;
assign equals_u22=equals_u22_a_signed==equals_u22_b_signed;
assign andOp_u29=equals_u21&equals_u22;
assign equals_u23_a_unsigned=port_2e0d86cd_;
assign equals_u23_b_unsigned=32'h20000;
assign equals_u23=equals_u23_a_unsigned==equals_u23_b_unsigned;
assign andOp_u30=andOp_u29&equals_u23;
assign andOp_u31=andOp_u30&port_70e1f405_;
assign equals_u24_a_unsigned=port_34f62b85_;
assign equals_u24_b_unsigned=16'h0;
assign equals_u24=equals_u24_a_unsigned==equals_u24_b_unsigned;
assign equals_u25_a_signed=port_6d2bfa2d_;
assign equals_u25_b_signed=16'h1ff;
assign equals_u25=equals_u25_a_signed==equals_u25_b_signed;
assign andOp_u32=equals_u24&equals_u25;
assign equals_u26_a_unsigned=port_2e0d86cd_;
assign equals_u26_b_unsigned=32'h20000;
assign equals_u26=equals_u26_a_unsigned==equals_u26_b_unsigned;
assign andOp_u33=andOp_u32&equals_u26;
assign not_u60=!port_70e1f405_;
assign andOp_u34=andOp_u33&not_u60;
assign lessThan_u17_a_unsigned=port_34f62b85_;
assign lessThan_u17_b_unsigned=16'hff;
assign lessThan_u17=lessThan_u17_a_unsigned<lessThan_u17_b_unsigned;
assign equals_u27_a_unsigned=port_2e0d86cd_;
assign equals_u27_b_unsigned=32'h20000;
assign equals_u27=equals_u27_a_unsigned==equals_u27_b_unsigned;
assign andOp_u35=lessThan_u17&equals_u27;
assign andOp_u36=andOp_u35&port_70e1f405_;
assign lessThan_u18_a_unsigned=port_34f62b85_;
assign lessThan_u18_b_unsigned=16'hff;
assign lessThan_u18=lessThan_u18_a_unsigned<lessThan_u18_b_unsigned;
assign equals_u28_a_unsigned=port_2e0d86cd_;
assign equals_u28_b_unsigned=32'h20000;
assign equals_u28=equals_u28_a_unsigned==equals_u28_b_unsigned;
assign andOp_u37=lessThan_u18&equals_u28;
assign not_u61=!port_70e1f405_;
assign andOp_u38=andOp_u37&not_u61;
assign equals_u29_a_unsigned=port_34f62b85_;
assign equals_u29_b_unsigned=16'hff;
assign equals_u29=equals_u29_a_unsigned==equals_u29_b_unsigned;
assign equals_u30_a_unsigned=port_2e0d86cd_;
assign equals_u30_b_unsigned=32'h20000;
assign equals_u30=equals_u30_a_unsigned==equals_u30_b_unsigned;
assign andOp_u39=equals_u29&equals_u30;
assign andOp_u40=andOp_u39&port_70e1f405_;
assign equals_u31_a_unsigned=port_34f62b85_;
assign equals_u31_b_unsigned=16'hff;
assign equals_u31=equals_u31_a_unsigned==equals_u31_b_unsigned;
assign equals_u32_a_unsigned=port_2e0d86cd_;
assign equals_u32_b_unsigned=32'h20000;
assign equals_u32=equals_u32_a_unsigned==equals_u32_b_unsigned;
assign andOp_u41=equals_u31&equals_u32;
assign not_u62=!port_70e1f405_;
assign andOp_u42=andOp_u41&not_u62;
assign equals_u33_a_signed={29'b0, port_42620ba7_};
assign equals_u33_b_signed=32'h0;
assign equals_u33=equals_u33_a_signed==equals_u33_b_signed;
assign and_u392_u0=and_u391_u0&not_u63_u0;
assign not_u63_u0=~equals_u33;
assign and_u393_u0=and_u391_u0&equals_u33;
assign andOp_u43=lessThan&port_6d3af1f9_;
assign not_u64_u0=~andOp_u43;
assign and_u394_u0=and_u401_u0&andOp_u43;
assign and_u395_u0=and_u401_u0&not_u64_u0;
assign simplePinWrite=and_u399_u0&{1{and_u399_u0}};
assign and_u396_u0=and_u400_u0&not_u65_u0;
assign not_u65_u0=~equals;
assign and_u397_u0=and_u400_u0&equals;
assign simplePinWrite_u74=and_u398_u0&{1{and_u398_u0}};
assign and_u398_u0=and_u397_u0&and_u400_u0;
assign and_u399_u0=and_u394_u0&and_u401_u0;
assign or_u86_u0=and_u399_u0|and_u398_u0;
assign mux_u28=(and_u399_u0)?3'h0:3'h1;
assign and_u400_u0=and_u395_u0&and_u401_u0;
assign and_u401_u0=and_u393_u0&and_u391_u0;
assign equals_u34_a_signed={29'b0, port_42620ba7_};
assign equals_u34_b_signed=32'h1;
assign equals_u34=equals_u34_a_signed==equals_u34_b_signed;
assign and_u402_u0=and_u391_u0&equals_u34;
assign not_u66_u0=~equals_u34;
assign and_u403_u0=and_u391_u0&not_u66_u0;
assign and_u404_u0=and_u413_u0&not_u67_u0;
assign not_u67_u0=~port_6d3af1f9_;
assign and_u405_u0=and_u413_u0&port_6d3af1f9_;
assign and_u406_u0=and_u411_u0&port_5e08959f_;
assign and_u407_u0=and_u411_u0&not_u68_u0;
assign not_u68_u0=~port_5e08959f_;
assign simplePinWrite_u75=and_u408_u0&{1{and_u408_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3a1f45fa_u0<=1'h0;
else reg_3a1f45fa_u0<=and_u408_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_75145b92_u0<=1'h0;
else reg_75145b92_u0<=reg_3a1f45fa_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_747e49b6_u0<=1'h0;
else reg_747e49b6_u0<=and_u409_u0;
end
assign and_u408_u0=and_u406_u0&and_u411_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_33c17034_u0<=1'h0;
else reg_33c17034_u0<=reg_75145b92_result_delayed_u0;
end
assign and_u409_u0=and_u407_u0&and_u411_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_33c17034_result_delayed_u0<=1'h0;
else reg_33c17034_result_delayed_u0<=reg_33c17034_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3a1f45fa_result_delayed_u0<=1'h0;
else reg_3a1f45fa_result_delayed_u0<=reg_3a1f45fa_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_75145b92_result_delayed_u0<=1'h0;
else reg_75145b92_result_delayed_u0<=reg_75145b92_u0;
end
assign or_u87_u0=reg_33c17034_result_delayed_u0|reg_747e49b6_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_66d1b020_u0<=1'h0;
else reg_66d1b020_u0<=and_u410_u0;
end
assign and_u410_u0=and_u404_u0&and_u413_u0;
assign or_u88_u0=or_u87_u0|reg_66d1b020_u0;
assign and_u411_u0=and_u405_u0&and_u413_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1b67eb07_u0<=1'h0;
else reg_1b67eb07_u0<=and_u412_u0;
end
assign and_u412_u0=and_u403_u0&and_u391_u0;
assign and_u413_u0=and_u402_u0&and_u391_u0;
assign or_u89_u0=or_u88_u0|reg_1b67eb07_u0;
assign equals_u35_a_signed={29'b0, port_42620ba7_};
assign equals_u35_b_signed=32'h2;
assign equals_u35=equals_u35_a_signed==equals_u35_b_signed;
assign and_u414_u0=and_u391_u0&not_u69_u0;
assign not_u69_u0=~equals_u35;
assign and_u415_u0=and_u391_u0&equals_u35;
assign andOp_u44=lessThan_u0&port_6d3af1f9_;
assign not_u70_u0=~andOp_u44;
assign and_u416_u0=and_u432_u0&andOp_u44;
assign and_u417_u0=and_u432_u0&not_u70_u0;
assign and_u418_u0=and_u430_u0&not_u71_u0;
assign not_u71_u0=~port_5e08959f_;
assign and_u419_u0=and_u430_u0&port_5e08959f_;
assign simplePinWrite_u76=and_u421_u0&{1{and_u421_u0}};
assign and_u420_u0=and_u418_u0&and_u430_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_179dcff8_u0<=1'h0;
else reg_179dcff8_u0<=reg_0322b1ca_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7d7c20fb_u0<=1'h0;
else reg_7d7c20fb_u0<=and_u421_u0;
end
assign and_u421_u0=and_u419_u0&and_u430_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0322b1ca_u0<=1'h0;
else reg_0322b1ca_u0<=reg_7d7c20fb_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_38422e0b_u0<=1'h0;
else reg_38422e0b_u0<=reg_179dcff8_result_delayed_u0;
end
assign or_u90_u0=and_delayed_u4|reg_38422e0b_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u4<=1'h0;
else and_delayed_u4<=and_u420_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7d7c20fb_result_delayed_u0<=1'h0;
else reg_7d7c20fb_result_delayed_u0<=reg_7d7c20fb_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_179dcff8_result_delayed_u0<=1'h0;
else reg_179dcff8_result_delayed_u0<=reg_179dcff8_u0;
end
assign andOp_u45=equals_u6&port_6d3af1f9_;
assign and_u422_u0=and_u431_u0&not_u72_u0;
assign not_u72_u0=~andOp_u45;
assign and_u423_u0=and_u431_u0&andOp_u45;
assign and_u424_u0=and_u429_u0&port_5e08959f_;
assign and_u425_u0=and_u429_u0&not_u73_u0;
assign not_u73_u0=~port_5e08959f_;
assign simplePinWrite_u77=and_u426_u0&{1{and_u426_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6f660aa7_u0<=1'h0;
else reg_6f660aa7_u0<=reg_115cba2e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1a2c6ea5_u0<=1'h0;
else reg_1a2c6ea5_u0<=and_u426_u0;
end
assign or_u91_u0=reg_6f660aa7_result_delayed_result_delayed_u0|reg_2e392276_u0;
assign and_u426_u0=and_u424_u0&and_u429_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6f660aa7_result_delayed_u0<=1'h0;
else reg_6f660aa7_result_delayed_u0<=reg_6f660aa7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2e392276_u0<=1'h0;
else reg_2e392276_u0<=and_u427_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_115cba2e_u0<=1'h0;
else reg_115cba2e_u0<=reg_1a2c6ea5_result_delayed_u0;
end
assign and_u427_u0=and_u425_u0&and_u429_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1a2c6ea5_result_delayed_u0<=1'h0;
else reg_1a2c6ea5_result_delayed_u0<=reg_1a2c6ea5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6f660aa7_result_delayed_result_delayed_u0<=1'h0;
else reg_6f660aa7_result_delayed_result_delayed_u0<=reg_6f660aa7_result_delayed_u0;
end
assign and_u428_u0=and_u422_u0&and_u431_u0;
assign and_u429_u0=and_u423_u0&and_u431_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u5_u0<=1'h0;
else and_delayed_u5_u0<=and_u428_u0;
end
assign or_u92_u0=and_delayed_u5_u0|or_u91_u0;
assign or_u93_u0=and_u421_u0|and_u426_u0;
assign mux_u29_u0=(and_u421_u0)?3'h2:3'h3;
assign and_u430_u0=and_u416_u0&and_u432_u0;
assign or_u94_u0=or_u92_u0|or_u90_u0;
assign and_u431_u0=and_u417_u0&and_u432_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3f285a69_u0<=1'h0;
else reg_3f285a69_u0<=and_u433_u0;
end
assign and_u432_u0=and_u415_u0&and_u391_u0;
assign and_u433_u0=and_u414_u0&and_u391_u0;
assign or_u95_u0=reg_3f285a69_u0|or_u94_u0;
assign equals_u36_a_signed={29'b0, port_42620ba7_};
assign equals_u36_b_signed=32'h3;
assign equals_u36=equals_u36_a_signed==equals_u36_b_signed;
assign not_u74_u0=~equals_u36;
assign and_u434_u0=and_u391_u0&equals_u36;
assign and_u435_u0=and_u391_u0&not_u74_u0;
assign andOp_u46=andOp_u1&port_6d3af1f9_;
assign and_u436_u0=and_u468_u0&not_u75_u0;
assign and_u437_u0=and_u468_u0&andOp_u46;
assign not_u75_u0=~andOp_u46;
assign and_u438_u0=and_u466_u0&port_5e08959f_;
assign not_u76_u0=~port_5e08959f_;
assign and_u439_u0=and_u466_u0&not_u76_u0;
assign simplePinWrite_u78=and_u441_u0&{1{and_u441_u0}};
assign or_u96_u0=reg_6a7d31d4_result_delayed_result_delayed_u0|and_delayed_u6_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4fb73053_u0<=1'h0;
else reg_4fb73053_u0<=and_u441_u0;
end
assign and_u440_u0=and_u439_u0&and_u466_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6a7d31d4_u0<=1'h0;
else reg_6a7d31d4_u0<=reg_63ede03c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u6_u0<=1'h0;
else and_delayed_u6_u0<=and_u440_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_63ede03c_u0<=1'h0;
else reg_63ede03c_u0<=reg_4fb73053_result_delayed_u0;
end
assign and_u441_u0=and_u438_u0&and_u466_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4fb73053_result_delayed_u0<=1'h0;
else reg_4fb73053_result_delayed_u0<=reg_4fb73053_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6a7d31d4_result_delayed_u0<=1'h0;
else reg_6a7d31d4_result_delayed_u0<=reg_6a7d31d4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6a7d31d4_result_delayed_result_delayed_u0<=1'h0;
else reg_6a7d31d4_result_delayed_result_delayed_u0<=reg_6a7d31d4_result_delayed_u0;
end
assign andOp_u47=andOp_u4&port_6d3af1f9_;
assign not_u77_u0=~andOp_u47;
assign and_u442_u0=and_u467_u0&andOp_u47;
assign and_u443_u0=and_u467_u0&not_u77_u0;
assign and_u444_u0=and_u465_u0&port_0cc0d92d_;
assign not_u78_u0=~port_0cc0d92d_;
assign and_u445_u0=and_u465_u0&not_u78_u0;
assign simplePinWrite_u79=and_u447_u0&{1{and_u447_u0}};
assign and_u446_u0=and_u445_u0&and_u465_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4dff0c7d_u0<=1'h0;
else reg_4dff0c7d_u0<=and_u447_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4dff0c7d_result_delayed_u0<=1'h0;
else reg_4dff0c7d_result_delayed_u0<=reg_4dff0c7d_u0;
end
assign and_u447_u0=and_u444_u0&and_u465_u0;
assign or_u97_u0=reg_4056b2dd_result_delayed_u0|and_delayed_u7_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4056b2dd_u0<=1'h0;
else reg_4056b2dd_u0<=reg_0da41b16_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0da41b16_u0<=1'h0;
else reg_0da41b16_u0<=reg_4dff0c7d_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4dff0c7d_result_delayed_result_delayed_u0<=1'h0;
else reg_4dff0c7d_result_delayed_result_delayed_u0<=reg_4dff0c7d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u7_u0<=1'h0;
else and_delayed_u7_u0<=and_u446_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4056b2dd_result_delayed_u0<=1'h0;
else reg_4056b2dd_result_delayed_u0<=reg_4056b2dd_u0;
end
assign not_u79_u0=~andOp_u7;
assign and_u448_u0=and_u464_u0&andOp_u7;
assign and_u449_u0=and_u464_u0&not_u79_u0;
assign not_u80_u0=~port_5e08959f_;
assign and_u450_u0=and_u463_u0&port_5e08959f_;
assign and_u451_u0=and_u463_u0&not_u80_u0;
assign simplePinWrite_u80=and_u452_u0&{1{and_u452_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_39b080d6_u0<=1'h0;
else reg_39b080d6_u0<=and_u453_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_54f4b899_u0<=1'h0;
else reg_54f4b899_u0<=and_u452_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_54f4b899_result_delayed_u0<=1'h0;
else reg_54f4b899_result_delayed_u0<=reg_54f4b899_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_66a4207d_u0<=1'h0;
else reg_66a4207d_u0<=reg_7c85adb8_u0;
end
assign and_u452_u0=and_u450_u0&and_u463_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7c85adb8_u0<=1'h0;
else reg_7c85adb8_u0<=reg_54f4b899_result_delayed_result_delayed_u0;
end
assign or_u98_u0=reg_39b080d6_u0|reg_66a4207d_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_54f4b899_result_delayed_result_delayed_u0<=1'h0;
else reg_54f4b899_result_delayed_result_delayed_u0<=reg_54f4b899_result_delayed_u0;
end
assign and_u453_u0=and_u451_u0&and_u463_u0;
assign and_u454_u0=and_u462_u0&andOp_u10;
assign and_u455_u0=and_u462_u0&not_u81_u0;
assign not_u81_u0=~andOp_u10;
assign and_u456_u0=and_u461_u0&not_u82_u0;
assign and_u457_u0=and_u461_u0&port_0cc0d92d_;
assign not_u82_u0=~port_0cc0d92d_;
assign simplePinWrite_u81=and_u459_u0&{1{and_u459_u0}};
assign and_u458_u0=and_u456_u0&and_u461_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_67690009_u0<=1'h0;
else reg_67690009_u0<=reg_2eb38cd6_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2eb38cd6_u0<=1'h0;
else reg_2eb38cd6_u0<=and_delayed_u9_u0;
end
assign or_u99_u0=and_delayed_u8_u0|reg_67690009_result_delayed_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u8_u0<=1'h0;
else and_delayed_u8_u0<=and_u458_u0;
end
assign and_u459_u0=and_u457_u0&and_u461_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2eb38cd6_result_delayed_u0<=1'h0;
else reg_2eb38cd6_result_delayed_u0<=reg_2eb38cd6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_67690009_result_delayed_u0<=1'h0;
else reg_67690009_result_delayed_u0<=reg_67690009_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u9_u0<=1'h0;
else and_delayed_u9_u0<=and_u459_u0;
end
assign and_u460_u0=and_u455_u0&and_u462_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u10_u0<=1'h0;
else and_delayed_u10_u0<=and_u460_u0;
end
assign or_u100_u0=or_u99_u0|and_delayed_u10_u0;
assign and_u461_u0=and_u454_u0&and_u462_u0;
assign or_u101_u0=or_u98_u0|or_u100_u0;
assign and_u462_u0=and_u449_u0&and_u464_u0;
assign and_u463_u0=and_u448_u0&and_u464_u0;
assign or_u102_u0=and_u452_u0|and_u459_u0;
assign and_u464_u0=and_u443_u0&and_u467_u0;
assign or_u103_u0=and_u447_u0|or_u102_u0;
assign or_u104_u0=or_u97_u0|or_u101_u0;
assign and_u465_u0=and_u442_u0&and_u467_u0;
assign or_u105_u0=or_u96_u0|or_u104_u0;
assign and_u466_u0=and_u437_u0&and_u468_u0;
assign and_u467_u0=and_u436_u0&and_u468_u0;
assign or_u106_u0=and_u441_u0|or_u103_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4e472843_u0<=1'h0;
else reg_4e472843_u0<=and_u469_u0;
end
assign and_u468_u0=and_u434_u0&and_u391_u0;
assign and_u469_u0=and_u435_u0&and_u391_u0;
assign or_u107_u0=or_u105_u0|reg_4e472843_u0;
assign equals_u37_a_signed={29'b0, port_42620ba7_};
assign equals_u37_b_signed=32'h4;
assign equals_u37=equals_u37_a_signed==equals_u37_b_signed;
assign and_u470_u0=and_u391_u0&equals_u37;
assign and_u471_u0=and_u391_u0&not_u83_u0;
assign not_u83_u0=~equals_u37;
assign andOp_u48=andOp_u13&port_6d3af1f9_;
assign and_u472_u0=and_u536_u0&not_u84_u0;
assign not_u84_u0=~andOp_u48;
assign and_u473_u0=and_u536_u0&andOp_u48;
assign not_u85_u0=~port_5e08959f_;
assign and_u474_u0=and_u534_u0&not_u85_u0;
assign and_u475_u0=and_u534_u0&port_5e08959f_;
assign simplePinWrite_u82=and_u476_u0&{1{and_u476_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6e3a0db9_u0<=1'h0;
else reg_6e3a0db9_u0<=reg_4d5434d2_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_43d57d30_u0<=1'h0;
else reg_43d57d30_u0<=and_u477_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4d5434d2_u0<=1'h0;
else reg_4d5434d2_u0<=reg_5bff6a34_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5bff6a34_u0<=1'h0;
else reg_5bff6a34_u0<=and_u476_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5bff6a34_result_delayed_u0<=1'h0;
else reg_5bff6a34_result_delayed_u0<=reg_5bff6a34_u0;
end
assign or_u108_u0=reg_6e3a0db9_u0|reg_43d57d30_u0;
assign and_u476_u0=and_u475_u0&and_u534_u0;
assign and_u477_u0=and_u474_u0&and_u534_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5bff6a34_result_delayed_result_delayed_u0<=1'h0;
else reg_5bff6a34_result_delayed_result_delayed_u0<=reg_5bff6a34_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4d5434d2_result_delayed_u0<=1'h0;
else reg_4d5434d2_result_delayed_u0<=reg_4d5434d2_u0;
end
assign andOp_u49=andOp_u16&port_6d3af1f9_;
assign and_u478_u0=and_u535_u0&not_u86_u0;
assign not_u86_u0=~andOp_u49;
assign and_u479_u0=and_u535_u0&andOp_u49;
assign not_u87_u0=~port_0cc0d92d_;
assign and_u480_u0=and_u533_u0&not_u87_u0;
assign and_u481_u0=and_u533_u0&port_0cc0d92d_;
assign simplePinWrite_u83=and_u483_u0&{1{and_u483_u0}};
assign or_u109_u0=reg_7b478222_u0|reg_48ed0ea7_result_delayed_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7b478222_u0<=1'h0;
else reg_7b478222_u0<=and_u482_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2e3fd957_u0<=1'h0;
else reg_2e3fd957_u0<=and_u483_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_48ed0ea7_u0<=1'h0;
else reg_48ed0ea7_u0<=reg_6b6f3e79_u0;
end
assign and_u482_u0=and_u480_u0&and_u533_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_48ed0ea7_result_delayed_u0<=1'h0;
else reg_48ed0ea7_result_delayed_u0<=reg_48ed0ea7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6b6f3e79_u0<=1'h0;
else reg_6b6f3e79_u0<=reg_2e3fd957_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2e3fd957_result_delayed_u0<=1'h0;
else reg_2e3fd957_result_delayed_u0<=reg_2e3fd957_u0;
end
assign and_u483_u0=and_u481_u0&and_u533_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2e3fd957_result_delayed_result_delayed_u0<=1'h0;
else reg_2e3fd957_result_delayed_result_delayed_u0<=reg_2e3fd957_result_delayed_u0;
end
assign not_u88_u0=~andOp_u18;
assign and_u484_u0=and_u532_u0&andOp_u18;
assign and_u485_u0=and_u532_u0&not_u88_u0;
assign not_u89_u0=~port_5e08959f_;
assign and_u486_u0=and_u531_u0&not_u89_u0;
assign and_u487_u0=and_u531_u0&port_5e08959f_;
assign simplePinWrite_u84=and_u489_u0&{1{and_u489_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6d9aed1d_u0<=1'h0;
else reg_6d9aed1d_u0<=reg_1decc03f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5afb3453_u0<=1'h0;
else reg_5afb3453_u0<=and_u488_u0;
end
assign and_u488_u0=and_u486_u0&and_u531_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1c6adbe7_u0<=1'h0;
else reg_1c6adbe7_u0<=reg_6d9aed1d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6d9aed1d_result_delayed_u0<=1'h0;
else reg_6d9aed1d_result_delayed_u0<=reg_6d9aed1d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1decc03f_u0<=1'h0;
else reg_1decc03f_u0<=and_u489_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1decc03f_result_delayed_u0<=1'h0;
else reg_1decc03f_result_delayed_u0<=reg_1decc03f_u0;
end
assign and_u489_u0=and_u487_u0&and_u531_u0;
assign or_u110_u0=reg_5afb3453_u0|reg_1c6adbe7_u0;
assign not_u90_u0=~andOp_u20;
assign and_u490_u0=and_u530_u0&andOp_u20;
assign and_u491_u0=and_u530_u0&not_u90_u0;
assign and_u492_u0=and_u528_u0&port_0cc0d92d_;
assign not_u91_u0=~port_0cc0d92d_;
assign and_u493_u0=and_u528_u0&not_u91_u0;
assign simplePinWrite_u85=and_u494_u0&{1{and_u494_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2b6f460f_u0<=1'h0;
else reg_2b6f460f_u0<=reg_4138b0a0_u0;
end
assign and_u494_u0=and_u492_u0&and_u528_u0;
assign and_u495_u0=and_u493_u0&and_u528_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2b6f460f_result_delayed_u0<=1'h0;
else reg_2b6f460f_result_delayed_u0<=reg_2b6f460f_u0;
end
assign or_u111_u0=and_delayed_u11_u0|reg_2b6f460f_result_delayed_result_delayed_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2b6f460f_result_delayed_result_delayed_u0<=1'h0;
else reg_2b6f460f_result_delayed_result_delayed_u0<=reg_2b6f460f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4138b0a0_u0<=1'h0;
else reg_4138b0a0_u0<=and_delayed_u12_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u11_u0<=1'h0;
else and_delayed_u11_u0<=and_u495_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u12_u0<=1'h0;
else and_delayed_u12_u0<=and_u494_u0;
end
assign andOp_u50=andOp_u22&port_6d3af1f9_;
assign and_u496_u0=and_u529_u0&andOp_u50;
assign not_u92_u0=~andOp_u50;
assign and_u497_u0=and_u529_u0&not_u92_u0;
assign and_u498_u0=and_u526_u0&not_u93_u0;
assign and_u499_u0=and_u526_u0&port_5e08959f_;
assign not_u93_u0=~port_5e08959f_;
assign simplePinWrite_u86=and_u501_u0&{1{and_u501_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5475b2b5_u0<=1'h0;
else reg_5475b2b5_u0<=and_u500_u0;
end
assign and_u500_u0=and_u498_u0&and_u526_u0;
assign and_u501_u0=and_u499_u0&and_u526_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7c3d02d5_u0<=1'h0;
else reg_7c3d02d5_u0<=and_delayed_u13_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7c3d02d5_result_delayed_u0<=1'h0;
else reg_7c3d02d5_result_delayed_u0<=reg_7c3d02d5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_424c04bc_u0<=1'h0;
else reg_424c04bc_u0<=reg_7c3d02d5_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_424c04bc_result_delayed_u0<=1'h0;
else reg_424c04bc_result_delayed_u0<=reg_424c04bc_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7c3d02d5_result_delayed_result_delayed_u0<=1'h0;
else reg_7c3d02d5_result_delayed_result_delayed_u0<=reg_7c3d02d5_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u13_u0<=1'h0;
else and_delayed_u13_u0<=and_u501_u0;
end
assign or_u112_u0=reg_424c04bc_result_delayed_u0|reg_5475b2b5_u0;
assign andOp_u51=andOp_u24&port_6d3af1f9_;
assign not_u94_u0=~andOp_u51;
assign and_u502_u0=and_u527_u0&andOp_u51;
assign and_u503_u0=and_u527_u0&not_u94_u0;
assign and_u504_u0=and_u524_u0&port_0cc0d92d_;
assign not_u95_u0=~port_0cc0d92d_;
assign and_u505_u0=and_u524_u0&not_u95_u0;
assign simplePinWrite_u87=and_u507_u0&{1{and_u507_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_71b65551_u0<=1'h0;
else reg_71b65551_u0<=reg_5557b19e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5557b19e_u0<=1'h0;
else reg_5557b19e_u0<=and_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_117d0bd6_u0<=1'h0;
else reg_117d0bd6_u0<=and_u506_u0;
end
assign or_u113_u0=reg_71b65551_result_delayed_u0|reg_117d0bd6_u0;
assign and_u506_u0=and_u505_u0&and_u524_u0;
assign and_u507_u0=and_u504_u0&and_u524_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u14_u0<=1'h0;
else and_delayed_u14_u0<=and_u507_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_result_delayed_u0<=1'h0;
else and_delayed_result_delayed_u0<=and_delayed_u14_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_71b65551_result_delayed_u0<=1'h0;
else reg_71b65551_result_delayed_u0<=reg_71b65551_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_result_delayed_result_delayed_u0<=1'h0;
else and_delayed_result_delayed_result_delayed_u0<=and_delayed_result_delayed_u0;
end
assign and_u508_u0=and_u525_u0&andOp_u26;
assign and_u509_u0=and_u525_u0&not_u96_u0;
assign not_u96_u0=~andOp_u26;
assign and_u510_u0=and_u523_u0&port_5e08959f_;
assign not_u97_u0=~port_5e08959f_;
assign and_u511_u0=and_u523_u0&not_u97_u0;
assign simplePinWrite_u88=and_u513_u0&{1{and_u513_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_04f3c4f4_u0<=1'h0;
else reg_04f3c4f4_u0<=reg_76e06d48_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_76e06d48_u0<=1'h0;
else reg_76e06d48_u0<=reg_7d698f03_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7d698f03_u0<=1'h0;
else reg_7d698f03_u0<=and_u513_u0;
end
assign and_u512_u0=and_u511_u0&and_u523_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7d698f03_result_delayed_u0<=1'h0;
else reg_7d698f03_result_delayed_u0<=reg_7d698f03_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u15_u0<=1'h0;
else and_delayed_u15_u0<=and_u512_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_04f3c4f4_result_delayed_u0<=1'h0;
else reg_04f3c4f4_result_delayed_u0<=reg_04f3c4f4_u0;
end
assign or_u114_u0=and_delayed_u15_u0|reg_04f3c4f4_result_delayed_u0;
assign and_u513_u0=and_u510_u0&and_u523_u0;
assign and_u514_u0=and_u522_u0&not_u98_u0;
assign not_u98_u0=~andOp_u28;
assign and_u515_u0=and_u522_u0&andOp_u28;
assign and_u516_u0=and_u521_u0&not_u99_u0;
assign and_u517_u0=and_u521_u0&port_0cc0d92d_;
assign not_u99_u0=~port_0cc0d92d_;
assign simplePinWrite_u89=and_u518_u0&{1{and_u518_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5b4fb5ce_u0<=1'h0;
else reg_5b4fb5ce_u0<=reg_52c1fee5_u0;
end
assign and_u518_u0=and_u517_u0&and_u521_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_52c1fee5_u0<=1'h0;
else reg_52c1fee5_u0<=reg_1ccb0e6e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1ccb0e6e_u0<=1'h0;
else reg_1ccb0e6e_u0<=and_delayed_u16_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u16_u0<=1'h0;
else and_delayed_u16_u0<=and_u518_u0;
end
assign or_u115_u0=reg_5b4fb5ce_result_delayed_u0|reg_26f8fd95_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_26f8fd95_u0<=1'h0;
else reg_26f8fd95_u0<=and_u519_u0;
end
assign and_u519_u0=and_u516_u0&and_u521_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5b4fb5ce_result_delayed_u0<=1'h0;
else reg_5b4fb5ce_result_delayed_u0<=reg_5b4fb5ce_u0;
end
assign and_u520_u0=and_u514_u0&and_u522_u0;
assign or_u116_u0=or_u115_u0|and_delayed_u17_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u17_u0<=1'h0;
else and_delayed_u17_u0<=and_u520_u0;
end
assign and_u521_u0=and_u515_u0&and_u522_u0;
assign and_u522_u0=and_u509_u0&and_u525_u0;
assign and_u523_u0=and_u508_u0&and_u525_u0;
assign or_u117_u0=or_u116_u0|or_u114_u0;
assign or_u118_u0=and_u513_u0|and_u518_u0;
assign or_u119_u0=or_u113_u0|or_u117_u0;
assign or_u120_u0=and_u507_u0|or_u118_u0;
assign and_u524_u0=and_u502_u0&and_u527_u0;
assign and_u525_u0=and_u503_u0&and_u527_u0;
assign and_u526_u0=and_u496_u0&and_u529_u0;
assign or_u121_u0=or_u112_u0|or_u119_u0;
assign or_u122_u0=and_u501_u0|or_u120_u0;
assign and_u527_u0=and_u497_u0&and_u529_u0;
assign mux_u30_u0=(and_u494_u0)?3'h4:3'h5;
assign or_u123_u0=and_u494_u0|or_u122_u0;
assign and_u528_u0=and_u490_u0&and_u530_u0;
assign or_u124_u0=or_u121_u0|or_u111_u0;
assign and_u529_u0=and_u491_u0&and_u530_u0;
assign and_u530_u0=and_u485_u0&and_u532_u0;
assign and_u531_u0=and_u484_u0&and_u532_u0;
assign or_u125_u0=and_u489_u0|or_u123_u0;
assign mux_u31_u0=(and_u489_u0)?3'h4:{2'b10, mux_u30_u0[0]};
assign or_u126_u0=or_u110_u0|or_u124_u0;
assign and_u532_u0=and_u478_u0&and_u535_u0;
assign and_u533_u0=and_u479_u0&and_u535_u0;
assign or_u127_u0=or_u126_u0|or_u109_u0;
assign or_u128_u0=and_u483_u0|or_u125_u0;
assign mux_u32_u0=(and_u483_u0)?3'h4:{2'b10, mux_u31_u0[0]};
assign and_u534_u0=and_u473_u0&and_u536_u0;
assign and_u535_u0=and_u472_u0&and_u536_u0;
assign or_u129_u0=and_u476_u0|or_u128_u0;
assign mux_u33_u0=(and_u476_u0)?3'h4:{2'b10, mux_u32_u0[0]};
assign or_u130_u0=or_u108_u0|or_u127_u0;
assign or_u131_u0=or_u130_u0|and_delayed_u18_u0;
assign and_u536_u0=and_u470_u0&and_u391_u0;
assign and_u537_u0=and_u471_u0&and_u391_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u18_u0<=1'h0;
else and_delayed_u18_u0<=and_u537_u0;
end
assign equals_u38_a_signed={29'b0, port_42620ba7_};
assign equals_u38_b_signed=32'h5;
assign equals_u38=equals_u38_a_signed==equals_u38_b_signed;
assign not_u100_u0=~equals_u38;
assign and_u538_u0=and_u391_u0&equals_u38;
assign and_u539_u0=and_u391_u0&not_u100_u0;
assign andOp_u52=andOp_u1&port_6d3af1f9_;
assign and_u540_u0=and_u588_u0&not_u101_u0;
assign not_u101_u0=~andOp_u52;
assign and_u541_u0=and_u588_u0&andOp_u52;
assign not_u102_u0=~port_5e08959f_;
assign and_u542_u0=and_u587_u0&port_5e08959f_;
assign and_u543_u0=and_u587_u0&not_u102_u0;
assign simplePinWrite_u90=and_u545_u0&{1{and_u545_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_60e797c7_u0<=1'h0;
else reg_60e797c7_u0<=reg_14bc455b_result_delayed_u0;
end
assign or_u132_u0=reg_60e797c7_u0|and_delayed_u19_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_14bc455b_u0<=1'h0;
else reg_14bc455b_u0<=reg_01c7fa9c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_14bc455b_result_delayed_u0<=1'h0;
else reg_14bc455b_result_delayed_u0<=reg_14bc455b_u0;
end
assign and_u544_u0=and_u543_u0&and_u587_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u19_u0<=1'h0;
else and_delayed_u19_u0<=and_u544_u0;
end
assign and_u545_u0=and_u542_u0&and_u587_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u20_u0<=1'h0;
else and_delayed_u20_u0<=and_u545_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01c7fa9c_u0<=1'h0;
else reg_01c7fa9c_u0<=and_delayed_result_delayed_u1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_result_delayed_u1_u0<=1'h0;
else and_delayed_result_delayed_u1_u0<=and_delayed_u20_u0;
end
assign andOp_u53=andOp_u4&port_6d3af1f9_;
assign and_u546_u0=and_u586_u0&not_u103_u0;
assign and_u547_u0=and_u586_u0&andOp_u53;
assign not_u103_u0=~andOp_u53;
assign and_u548_u0=and_u585_u0&port_0cc0d92d_;
assign and_u549_u0=and_u585_u0&not_u104_u0;
assign not_u104_u0=~port_0cc0d92d_;
assign simplePinWrite_u91=and_u550_u0&{1{and_u550_u0}};
assign and_u550_u0=and_u548_u0&and_u585_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7b1e075a_u0<=1'h0;
else reg_7b1e075a_u0<=and_delayed_u21_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_37e60342_u0<=1'h0;
else reg_37e60342_u0<=reg_7b1e075a_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0834cf70_u0<=1'h0;
else reg_0834cf70_u0<=and_u551_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_37e60342_result_delayed_u0<=1'h0;
else reg_37e60342_result_delayed_u0<=reg_37e60342_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7b1e075a_result_delayed_u0<=1'h0;
else reg_7b1e075a_result_delayed_u0<=reg_7b1e075a_u0;
end
assign and_u551_u0=and_u549_u0&and_u585_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7b1e075a_result_delayed_result_delayed_u0<=1'h0;
else reg_7b1e075a_result_delayed_result_delayed_u0<=reg_7b1e075a_result_delayed_u0;
end
assign or_u133_u0=reg_37e60342_result_delayed_u0|reg_0834cf70_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u21_u0<=1'h0;
else and_delayed_u21_u0<=and_u550_u0;
end
assign and_u552_u0=and_u584_u0&andOp_u7;
assign and_u553_u0=and_u584_u0&not_u105_u0;
assign not_u105_u0=~andOp_u7;
assign and_u554_u0=and_u582_u0&not_u106_u0;
assign and_u555_u0=and_u582_u0&port_5e08959f_;
assign not_u106_u0=~port_5e08959f_;
assign simplePinWrite_u92=and_u556_u0&{1{and_u556_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2b889e88_u0<=1'h0;
else reg_2b889e88_u0<=and_u556_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3fd6f110_u0<=1'h0;
else reg_3fd6f110_u0<=reg_2b889e88_result_delayed_u0;
end
assign and_u556_u0=and_u555_u0&and_u582_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_33af66c3_u0<=1'h0;
else reg_33af66c3_u0<=reg_3fd6f110_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2b889e88_result_delayed_u0<=1'h0;
else reg_2b889e88_result_delayed_u0<=reg_2b889e88_u0;
end
assign and_u557_u0=and_u554_u0&and_u582_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u22_u0<=1'h0;
else and_delayed_u22_u0<=and_u557_u0;
end
assign or_u134_u0=reg_33af66c3_u0|and_delayed_u22_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3fd6f110_result_delayed_u0<=1'h0;
else reg_3fd6f110_result_delayed_u0<=reg_3fd6f110_u0;
end
assign not_u107_u0=~andOp_u10;
assign and_u558_u0=and_u583_u0&not_u107_u0;
assign and_u559_u0=and_u583_u0&andOp_u10;
assign and_u560_u0=and_u580_u0&not_u108_u0;
assign and_u561_u0=and_u580_u0&port_0cc0d92d_;
assign not_u108_u0=~port_0cc0d92d_;
assign simplePinWrite_u93=and_u563_u0&{1{and_u563_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_49ed7469_u0<=1'h0;
else reg_49ed7469_u0<=and_u563_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_575d09b8_u0<=1'h0;
else reg_575d09b8_u0<=reg_6efc1130_u0;
end
assign and_u562_u0=and_u560_u0&and_u580_u0;
assign and_u563_u0=and_u561_u0&and_u580_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6efc1130_u0<=1'h0;
else reg_6efc1130_u0<=reg_49ed7469_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_49ed7469_result_delayed_u0<=1'h0;
else reg_49ed7469_result_delayed_u0<=reg_49ed7469_u0;
end
assign or_u135_u0=reg_575d09b8_u0|and_delayed_u23_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_49ed7469_result_delayed_result_delayed_u0<=1'h0;
else reg_49ed7469_result_delayed_result_delayed_u0<=reg_49ed7469_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u23_u0<=1'h0;
else and_delayed_u23_u0<=and_u562_u0;
end
assign and_u564_u0=and_u581_u0&andOp_u31;
assign not_u109_u0=~andOp_u31;
assign and_u565_u0=and_u581_u0&not_u109_u0;
assign and_u566_u0=and_u578_u0&not_u110_u0;
assign and_u567_u0=and_u578_u0&port_5e08959f_;
assign not_u110_u0=~port_5e08959f_;
assign simplePinWrite_u94=and_u569_u0&{1{and_u569_u0}};
assign and_u568_u0=and_u566_u0&and_u578_u0;
assign and_u569_u0=and_u567_u0&and_u578_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u24_u0<=1'h0;
else and_delayed_u24_u0<=and_u568_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1723f867_u0<=1'h0;
else reg_1723f867_u0<=reg_11292ccc_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_11292ccc_u0<=1'h0;
else reg_11292ccc_u0<=and_delayed_u25_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_11292ccc_result_delayed_u0<=1'h0;
else reg_11292ccc_result_delayed_u0<=reg_11292ccc_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u25_u0<=1'h0;
else and_delayed_u25_u0<=and_u569_u0;
end
assign or_u136_u0=reg_1723f867_u0|and_delayed_u24_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_11292ccc_result_delayed_result_delayed_u0<=1'h0;
else reg_11292ccc_result_delayed_result_delayed_u0<=reg_11292ccc_result_delayed_u0;
end
assign and_u570_u0=and_u579_u0&not_u111_u0;
assign and_u571_u0=and_u579_u0&andOp_u34;
assign not_u111_u0=~andOp_u34;
assign not_u112_u0=~port_0cc0d92d_;
assign and_u572_u0=and_u576_u0&port_0cc0d92d_;
assign and_u573_u0=and_u576_u0&not_u112_u0;
assign simplePinWrite_u95=and_u574_u0&{1{and_u574_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_64e07a44_u0<=1'h0;
else reg_64e07a44_u0<=and_u575_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_23dba81c_u0<=1'h0;
else reg_23dba81c_u0<=and_u574_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_23dba81c_result_delayed_u0<=1'h0;
else reg_23dba81c_result_delayed_u0<=reg_23dba81c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_15bcd7f0_u0<=1'h0;
else reg_15bcd7f0_u0<=reg_53451f0b_u0;
end
assign and_u574_u0=and_u572_u0&and_u576_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_53451f0b_u0<=1'h0;
else reg_53451f0b_u0<=reg_23dba81c_result_delayed_result_delayed_u0;
end
assign and_u575_u0=and_u573_u0&and_u576_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_23dba81c_result_delayed_result_delayed_u0<=1'h0;
else reg_23dba81c_result_delayed_result_delayed_u0<=reg_23dba81c_result_delayed_u0;
end
assign or_u137_u0=reg_15bcd7f0_u0|reg_64e07a44_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_106be70b_u0<=1'h0;
else reg_106be70b_u0<=and_u577_u0;
end
assign and_u576_u0=and_u571_u0&and_u579_u0;
assign or_u138_u0=or_u137_u0|reg_106be70b_u0;
assign and_u577_u0=and_u570_u0&and_u579_u0;
assign or_u139_u0=and_u569_u0|and_u574_u0;
assign and_u578_u0=and_u564_u0&and_u581_u0;
assign and_u579_u0=and_u565_u0&and_u581_u0;
assign or_u140_u0=or_u138_u0|or_u136_u0;
assign and_u580_u0=and_u559_u0&and_u583_u0;
assign and_u581_u0=and_u558_u0&and_u583_u0;
assign or_u141_u0=and_u563_u0|or_u139_u0;
assign mux_u34_u0=(and_u563_u0)?3'h4:3'h6;
assign or_u142_u0=or_u140_u0|or_u135_u0;
assign and_u582_u0=and_u552_u0&and_u584_u0;
assign and_u583_u0=and_u553_u0&and_u584_u0;
assign mux_u35_u0=(and_u556_u0)?3'h4:{1'b1, mux_u34_u0[1], 1'b0};
assign or_u143_u0=and_u556_u0|or_u141_u0;
assign or_u144_u0=or_u134_u0|or_u142_u0;
assign and_u584_u0=and_u546_u0&and_u586_u0;
assign and_u585_u0=and_u547_u0&and_u586_u0;
assign mux_u36_u0=(and_u550_u0)?3'h4:{1'b1, mux_u35_u0[1], 1'b0};
assign or_u145_u0=and_u550_u0|or_u143_u0;
assign or_u146_u0=or_u133_u0|or_u144_u0;
assign and_u586_u0=and_u540_u0&and_u588_u0;
assign or_u147_u0=and_u545_u0|or_u145_u0;
assign mux_u37_u0=(and_u545_u0)?3'h4:{1'b1, mux_u36_u0[1], 1'b0};
assign and_u587_u0=and_u541_u0&and_u588_u0;
assign or_u148_u0=or_u146_u0|or_u132_u0;
assign or_u149_u0=reg_1032f60e_u0|or_u148_u0;
assign and_u588_u0=and_u538_u0&and_u391_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1032f60e_u0<=1'h0;
else reg_1032f60e_u0<=and_u589_u0;
end
assign and_u589_u0=and_u539_u0&and_u391_u0;
assign equals_u39_a_signed={29'b0, port_42620ba7_};
assign equals_u39_b_signed=32'h6;
assign equals_u39=equals_u39_a_signed==equals_u39_b_signed;
assign and_u590_u0=and_u391_u0&equals_u39;
assign and_u591_u0=and_u391_u0&not_u113_u0;
assign not_u113_u0=~equals_u39;
assign and_u592_u0=and_u624_u0&andOp_u36;
assign not_u114_u0=~andOp_u36;
assign and_u593_u0=and_u624_u0&not_u114_u0;
assign and_u594_u0=and_u622_u0&port_5e08959f_;
assign and_u595_u0=and_u622_u0&not_u115_u0;
assign not_u115_u0=~port_5e08959f_;
assign simplePinWrite_u96=and_u597_u0&{1{and_u597_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_631bc458_u0<=1'h0;
else reg_631bc458_u0<=reg_789509d9_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_67355df6_u0<=1'h0;
else reg_67355df6_u0<=reg_631bc458_result_delayed_u0;
end
assign or_u150_u0=reg_67355df6_u0|reg_07f5313f_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_07f5313f_u0<=1'h0;
else reg_07f5313f_u0<=and_u596_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_789509d9_u0<=1'h0;
else reg_789509d9_u0<=and_u597_u0;
end
assign and_u596_u0=and_u595_u0&and_u622_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_631bc458_result_delayed_u0<=1'h0;
else reg_631bc458_result_delayed_u0<=reg_631bc458_u0;
end
assign and_u597_u0=and_u594_u0&and_u622_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_789509d9_result_delayed_u0<=1'h0;
else reg_789509d9_result_delayed_u0<=reg_789509d9_u0;
end
assign not_u116_u0=~andOp_u38;
assign and_u598_u0=and_u623_u0&andOp_u38;
assign and_u599_u0=and_u623_u0&not_u116_u0;
assign and_u600_u0=and_u621_u0&port_0cc0d92d_;
assign and_u601_u0=and_u621_u0&not_u117_u0;
assign not_u117_u0=~port_0cc0d92d_;
assign simplePinWrite_u97=and_u603_u0&{1{and_u603_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_45853e06_u0<=1'h0;
else reg_45853e06_u0<=reg_00fcf046_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_45853e06_result_delayed_u0<=1'h0;
else reg_45853e06_result_delayed_u0<=reg_45853e06_u0;
end
assign and_u602_u0=and_u601_u0&and_u621_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00fcf046_u0<=1'h0;
else reg_00fcf046_u0<=and_delayed_u26_u0;
end
assign or_u151_u0=reg_45853e06_result_delayed_result_delayed_u0|and_delayed_u27_u0;
assign and_u603_u0=and_u600_u0&and_u621_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u26_u0<=1'h0;
else and_delayed_u26_u0<=and_u603_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u27_u0<=1'h0;
else and_delayed_u27_u0<=and_u602_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_45853e06_result_delayed_result_delayed_u0<=1'h0;
else reg_45853e06_result_delayed_result_delayed_u0<=reg_45853e06_result_delayed_u0;
end
assign and_u604_u0=and_u620_u0&andOp_u40;
assign not_u118_u0=~andOp_u40;
assign and_u605_u0=and_u620_u0&not_u118_u0;
assign and_u606_u0=and_u619_u0&not_u119_u0;
assign not_u119_u0=~port_5e08959f_;
assign and_u607_u0=and_u619_u0&port_5e08959f_;
assign simplePinWrite_u98=and_u609_u0&{1{and_u609_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4b138e52_u0<=1'h0;
else reg_4b138e52_u0<=and_u609_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6bcd16e4_u0<=1'h0;
else reg_6bcd16e4_u0<=reg_36c01350_result_delayed_u0;
end
assign and_u608_u0=and_u606_u0&and_u619_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_36c01350_u0<=1'h0;
else reg_36c01350_u0<=reg_4b138e52_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_36c01350_result_delayed_u0<=1'h0;
else reg_36c01350_result_delayed_u0<=reg_36c01350_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u28_u0<=1'h0;
else and_delayed_u28_u0<=and_u608_u0;
end
assign and_u609_u0=and_u607_u0&and_u619_u0;
assign or_u152_u0=and_delayed_u28_u0|reg_6bcd16e4_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4b138e52_result_delayed_u0<=1'h0;
else reg_4b138e52_result_delayed_u0<=reg_4b138e52_u0;
end
assign and_u610_u0=and_u618_u0&not_u120_u0;
assign not_u120_u0=~andOp_u42;
assign and_u611_u0=and_u618_u0&andOp_u42;
assign and_u612_u0=and_u616_u0&not_u121_u0;
assign and_u613_u0=and_u616_u0&port_0cc0d92d_;
assign not_u121_u0=~port_0cc0d92d_;
assign simplePinWrite_u99=and_u614_u0&{1{and_u614_u0}};
assign and_u614_u0=and_u613_u0&and_u616_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u29_u0<=1'h0;
else and_delayed_u29_u0<=and_u614_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_result_delayed_u2_u0<=1'h0;
else and_delayed_result_delayed_u2_u0<=and_delayed_u29_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_265a004b_u0<=1'h0;
else reg_265a004b_u0<=and_delayed_result_delayed_result_delayed_u1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_265a004b_result_delayed_u0<=1'h0;
else reg_265a004b_result_delayed_u0<=reg_265a004b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_60ff05ab_u0<=1'h0;
else reg_60ff05ab_u0<=and_u615_u0;
end
assign and_u615_u0=and_u612_u0&and_u616_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_result_delayed_result_delayed_u1_u0<=1'h0;
else and_delayed_result_delayed_result_delayed_u1_u0<=and_delayed_result_delayed_u2_u0;
end
assign or_u153_u0=reg_265a004b_result_delayed_u0|reg_60ff05ab_u0;
assign and_u616_u0=and_u611_u0&and_u618_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_20083bde_u0<=1'h0;
else reg_20083bde_u0<=and_u617_u0;
end
assign and_u617_u0=and_u610_u0&and_u618_u0;
assign or_u154_u0=or_u153_u0|reg_20083bde_u0;
assign and_u618_u0=and_u605_u0&and_u620_u0;
assign or_u155_u0=and_u609_u0|and_u614_u0;
assign and_u619_u0=and_u604_u0&and_u620_u0;
assign or_u156_u0=or_u152_u0|or_u154_u0;
assign and_u620_u0=and_u599_u0&and_u623_u0;
assign or_u157_u0=or_u156_u0|or_u151_u0;
assign and_u621_u0=and_u598_u0&and_u623_u0;
assign or_u158_u0=and_u603_u0|or_u155_u0;
assign mux_u38_u0=(and_u603_u0)?3'h6:3'h0;
assign or_u159_u0=or_u157_u0|or_u150_u0;
assign and_u622_u0=and_u592_u0&and_u624_u0;
assign or_u160_u0=and_u597_u0|or_u158_u0;
assign mux_u39_u0=(and_u597_u0)?3'h6:{mux_u38_u0[1], mux_u38_u0[1], 1'b0};
assign and_u623_u0=and_u593_u0&and_u624_u0;
assign and_u624_u0=and_u590_u0&and_u391_u0;
assign and_u625_u0=and_u591_u0&and_u391_u0;
assign or_u161_u0=or_u159_u0|and_delayed_u30_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u30_u0<=1'h0;
else and_delayed_u30_u0<=and_u625_u0;
end
assign midLeft2_go_merge=simplePinWrite_u79|simplePinWrite_u91;
assign midLeft1_go_merge=simplePinWrite_u78|simplePinWrite_u90;
assign midLeftNoConsume2_go_merge=simplePinWrite_u81|simplePinWrite_u93;
assign midLeftNoConsume1_go_merge=simplePinWrite_u80|simplePinWrite_u92;
assign scoreboard_45f1cb9d_and=scoreboard_45f1cb9d_resOr0&scoreboard_45f1cb9d_resOr1&scoreboard_45f1cb9d_resOr2&scoreboard_45f1cb9d_resOr3&scoreboard_45f1cb9d_resOr4&scoreboard_45f1cb9d_resOr5;
always @(posedge CLK)
begin
if (bus_384ef3c0_)
scoreboard_45f1cb9d_reg0<=1'h0;
else if (or_u89_u0)
scoreboard_45f1cb9d_reg0<=1'h1;
else scoreboard_45f1cb9d_reg0<=scoreboard_45f1cb9d_reg0;
end
assign scoreboard_45f1cb9d_resOr3=or_u131_u0|scoreboard_45f1cb9d_reg3;
assign bus_384ef3c0_=scoreboard_45f1cb9d_and|RESET;
assign scoreboard_45f1cb9d_resOr4=or_u95_u0|scoreboard_45f1cb9d_reg4;
assign scoreboard_45f1cb9d_resOr0=or_u89_u0|scoreboard_45f1cb9d_reg0;
always @(posedge CLK)
begin
if (bus_384ef3c0_)
scoreboard_45f1cb9d_reg1<=1'h0;
else if (or_u107_u0)
scoreboard_45f1cb9d_reg1<=1'h1;
else scoreboard_45f1cb9d_reg1<=scoreboard_45f1cb9d_reg1;
end
always @(posedge CLK)
begin
if (bus_384ef3c0_)
scoreboard_45f1cb9d_reg5<=1'h0;
else if (or_u161_u0)
scoreboard_45f1cb9d_reg5<=1'h1;
else scoreboard_45f1cb9d_reg5<=scoreboard_45f1cb9d_reg5;
end
always @(posedge CLK)
begin
if (bus_384ef3c0_)
scoreboard_45f1cb9d_reg3<=1'h0;
else if (or_u131_u0)
scoreboard_45f1cb9d_reg3<=1'h1;
else scoreboard_45f1cb9d_reg3<=scoreboard_45f1cb9d_reg3;
end
assign scoreboard_45f1cb9d_resOr2=or_u149_u0|scoreboard_45f1cb9d_reg2;
always @(posedge CLK)
begin
if (bus_384ef3c0_)
scoreboard_45f1cb9d_reg4<=1'h0;
else if (or_u95_u0)
scoreboard_45f1cb9d_reg4<=1'h1;
else scoreboard_45f1cb9d_reg4<=scoreboard_45f1cb9d_reg4;
end
assign scoreboard_45f1cb9d_resOr1=or_u107_u0|scoreboard_45f1cb9d_reg1;
always @(posedge CLK)
begin
if (bus_384ef3c0_)
scoreboard_45f1cb9d_reg2<=1'h0;
else if (or_u149_u0)
scoreboard_45f1cb9d_reg2<=1'h1;
else scoreboard_45f1cb9d_reg2<=scoreboard_45f1cb9d_reg2;
end
assign scoreboard_45f1cb9d_resOr5=or_u161_u0|scoreboard_45f1cb9d_reg5;
assign mux_u40_u0=({3{or_u86_u0}}&{2'b0, mux_u28[0]})|({3{and_u408_u0}}&3'h2)|({3{or_u93_u0}}&{2'b1, mux_u29_u0[0]})|({3{or_u106_u0}}&3'h4)|({3{or_u129_u0}}&{2'b10, mux_u33_u0[0]})|({3{or_u147_u0}}&{1'b1, mux_u37_u0[1], 1'b0})|({3{or_u160_u0}}&{mux_u39_u0[1], mux_u39_u0[1], 1'b0});
assign or_u162_u0=or_u86_u0|and_u408_u0|or_u93_u0|or_u106_u0|or_u129_u0|or_u147_u0|or_u160_u0;
assign or_u163_u0=scoreboard_45f1cb9d_and|reg_45547147_result_delayed_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_45547147_u0<=1'h0;
else reg_45547147_u0<=GO;
end
assign mux_u41_u0=(GO)?3'h0:mux_u40_u0;
assign or_u164_u0=GO|or_u162_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_45547147_result_delayed_u0<=1'h0;
else reg_45547147_result_delayed_u0<=reg_45547147_u0;
end
assign RESULT=or_u164_u0;
assign RESULT_u320=mux_u41_u0;
assign RESULT_u321=midLeft1_go_merge;
assign RESULT_u322=simplePinWrite_u96;
assign RESULT_u323=simplePinWrite_u85;
assign RESULT_u324=simplePinWrite_u76;
assign RESULT_u325=simplePinWrite_u89;
assign RESULT_u326=simplePinWrite_u84;
assign RESULT_u327=simplePinWrite_u94;
assign RESULT_u328=simplePinWrite_u77;
assign RESULT_u329=midLeftNoConsume2_go_merge;
assign RESULT_u330=simplePinWrite_u95;
assign RESULT_u331=simplePinWrite_u99;
assign RESULT_u332=simplePinWrite_u83;
assign RESULT_u333=simplePinWrite_u97;
assign RESULT_u334=simplePinWrite_u82;
assign RESULT_u335=simplePinWrite_u88;
assign RESULT_u336=simplePinWrite_u98;
assign RESULT_u337=midLeft2_go_merge;
assign RESULT_u338=simplePinWrite;
assign RESULT_u339=midLeftNoConsume1_go_merge;
assign RESULT_u340=simplePinWrite_u87;
assign RESULT_u341=simplePinWrite_u86;
assign RESULT_u342=simplePinWrite_u75;
assign RESULT_u343=simplePinWrite_u74;
assign DONE=1'h0;
endmodule



module LL1_H_iunzipFilter2D_midRightNoConsume1(CLK, RESET, GO, port_5a871a00_, port_41319ec4_, port_462e5940_, port_7baa5f0a_, RESULT, RESULT_u344, RESULT_u345, RESULT_u346, RESULT_u347, RESULT_u348, RESULT_u349, RESULT_u350, RESULT_u351, RESULT_u352, RESULT_u353, RESULT_u354, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_5a871a00_;
input		port_41319ec4_;
input		port_462e5940_;
input	[15:0]	port_7baa5f0a_;
output		RESULT;
output	[15:0]	RESULT_u344;
output		RESULT_u345;
output	[15:0]	RESULT_u346;
output		RESULT_u347;
output		RESULT_u348;
output		RESULT_u349;
output	[31:0]	RESULT_u350;
output	[2:0]	RESULT_u351;
output	[15:0]	RESULT_u352;
output		RESULT_u353;
output	[15:0]	RESULT_u354;
output		DONE;
reg		done_cache_u38=1'h0;
wire		and_u627_u0;
wire		or_u165_u0;
wire		and_u632_u0;
wire		or_u166_u0;
reg		done_cache_u39_u0=1'h0;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_04ae8e2d_instance_RESULT;
wire	[15:0]	add;
wire		not_u123;
wire	[15:0]	simplePinWrite;
wire	[15:0]	simplePinWrite_u100;
wire		simplePinWrite_u101;
reg	[15:0]	syncEnable_u28=16'h0;
reg		reg_5cac2cfe_u0=1'h0;
reg		reg_24e2c079_u0=1'h0;
reg		reg_3b977622_u0=1'h0;
reg		reg_1a5485ed_u0=1'h0;
wire		or_u167_u0;
reg		reg_3b977622_result_delayed_u0=1'h0;
always @(posedge CLK or posedge GO or posedge or_u165_u0)
begin
if (or_u165_u0)
done_cache_u38<=1'h0;
else if (GO)
done_cache_u38<=1'h1;
else done_cache_u38<=done_cache_u38;
end
assign and_u627_u0=done_cache_u38&port_462e5940_;
assign or_u165_u0=and_u627_u0|RESET;
assign and_u632_u0=done_cache_u39_u0&port_462e5940_;
assign or_u166_u0=and_u632_u0|RESET;
always @(posedge CLK or posedge reg_3b977622_result_delayed_u0 or posedge or_u166_u0)
begin
if (or_u166_u0)
done_cache_u39_u0<=1'h0;
else if (reg_3b977622_result_delayed_u0)
done_cache_u39_u0<=1'h1;
else done_cache_u39_u0<=done_cache_u39_u0;
end
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_04ae8e2d_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_04ae8e2d_instance(.GO(reg_1a5485ed_u0), 
  .port_04d747de_(syncEnable_u28), .port_50018aab_(port_7baa5f0a_), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_04ae8e2d_instance_RESULT));
assign add=port_5a871a00_+16'h1;
assign not_u123=!port_41319ec4_;
assign simplePinWrite=16'h1&{16{1'h1}};
assign simplePinWrite_u100=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_04ae8e2d_instance_RESULT&{16{reg_1a5485ed_u0}};
assign simplePinWrite_u101=reg_1a5485ed_u0&{1{reg_1a5485ed_u0}};
always @(posedge CLK)
begin
if (reg_3b977622_u0)
syncEnable_u28<=port_7baa5f0a_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5cac2cfe_u0<=1'h0;
else reg_5cac2cfe_u0<=reg_24e2c079_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_24e2c079_u0<=1'h0;
else reg_24e2c079_u0<=reg_1a5485ed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3b977622_u0<=1'h0;
else reg_3b977622_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1a5485ed_u0<=1'h0;
else reg_1a5485ed_u0<=reg_3b977622_result_delayed_u0;
end
assign or_u167_u0=GO|reg_3b977622_result_delayed_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3b977622_result_delayed_u0<=1'h0;
else reg_3b977622_result_delayed_u0<=reg_3b977622_u0;
end
assign RESULT=GO;
assign RESULT_u344=add;
assign RESULT_u345=GO;
assign RESULT_u346=16'h0;
assign RESULT_u347=GO;
assign RESULT_u348=not_u123;
assign RESULT_u349=or_u167_u0;
assign RESULT_u350=32'h0;
assign RESULT_u351=3'h1;
assign RESULT_u352=simplePinWrite;
assign RESULT_u353=simplePinWrite_u101;
assign RESULT_u354=simplePinWrite_u100;
assign DONE=reg_5cac2cfe_u0;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_04ae8e2d_(GO, port_04d747de_, port_50018aab_, RESULT);
input		GO;
input	[15:0]	port_04d747de_;
input	[15:0]	port_50018aab_;
output	[15:0]	RESULT;
wire	[16:0]	add;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_3f570b28_instance_RESULT;
assign add={port_04d747de_[15], port_04d747de_}+{port_50018aab_[15], port_50018aab_};
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_3f570b28_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_3f570b28_instance(.GO(GO), 
  .port_3fbd9c0b_({add[16], add[16:2]}), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_3f570b28_instance_RESULT));
assign RESULT=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_3f570b28_instance_RESULT;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_3f570b28_(GO, port_3fbd9c0b_, RESULT);
input		GO;
input	[15:0]	port_3fbd9c0b_;
output	[15:0]	RESULT;
wire		greaterThan;
wire signed	[15:0]	greaterThan_b_signed;
wire signed	[15:0]	greaterThan_a_signed;
wire		and_u636_u0;
wire		and_u637_u0;
wire		not_u122_u0;
wire		and_u638_u0;
wire	[15:0]	mux_u42;
wire		and_u639_u0;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_3fbd9c0b_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign and_u636_u0=GO&greaterThan;
assign and_u637_u0=GO&not_u122_u0;
assign not_u122_u0=~greaterThan;
assign and_u638_u0=and_u636_u0&GO;
assign mux_u42=(and_u638_u0)?16'h0:port_3fbd9c0b_;
assign and_u639_u0=and_u637_u0&GO;
assign RESULT=mux_u42;
endmodule



module LL1_H_iunzipFilter2D_midRight1(CLK, RESET, GO, port_5330dddc_, port_0e198730_, port_55a91fbd_, port_4d6b8630_, port_610b7aeb_, port_0ba14e5d_, port_58e85b4e_, RESULT, RESULT_u355, RESULT_u356, RESULT_u357, RESULT_u358, RESULT_u359, RESULT_u360, RESULT_u361, RESULT_u362, RESULT_u363, RESULT_u364, RESULT_u365, RESULT_u366, RESULT_u367, RESULT_u368, RESULT_u369, RESULT_u370, RESULT_u371, RESULT_u372, RESULT_u373, RESULT_u374, DONE);
input		CLK;
input		RESET;
input		GO;
input	[31:0]	port_5330dddc_;
input	[15:0]	port_0e198730_;
input		port_55a91fbd_;
input		port_4d6b8630_;
input	[15:0]	port_610b7aeb_;
input		port_0ba14e5d_;
input	[15:0]	port_58e85b4e_;
output		RESULT;
output	[15:0]	RESULT_u355;
output		RESULT_u356;
output	[31:0]	RESULT_u357;
output		RESULT_u358;
output	[15:0]	RESULT_u359;
output		RESULT_u360;
output	[15:0]	RESULT_u361;
output		RESULT_u362;
output		RESULT_u363;
output		RESULT_u364;
output	[31:0]	RESULT_u365;
output	[2:0]	RESULT_u366;
output		RESULT_u367;
output	[31:0]	RESULT_u368;
output	[15:0]	RESULT_u369;
output	[2:0]	RESULT_u370;
output		RESULT_u371;
output	[15:0]	RESULT_u372;
output		RESULT_u373;
output	[15:0]	RESULT_u374;
output		DONE;
wire		simplePinWrite;
wire		and_u641_u0;
wire		or_u168_u0;
reg		done_cache_u40=1'h0;
wire		and_u646_u0;
reg		done_cache_u41_u0=1'h0;
wire		or_u169_u0;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_7779df0d_instance_RESULT;
reg		reg_663425d2_u0=1'h0;
wire		and_u655_u0;
wire		or_u170_u0;
wire	[31:0]	add;
wire	[15:0]	add_u11;
wire		not_u125;
wire		simplePinWrite_u102;
wire	[15:0]	simplePinWrite_u103;
wire	[15:0]	simplePinWrite_u104;
reg		reg_7fa5a9ca_u0=1'h0;
wire		or_u171_u0;
reg		reg_6857eec0_u0=1'h0;
reg		reg_644a10e2_u0=1'h0;
reg		reg_5a7b2b71_u0=1'h0;
reg		reg_644a10e2_result_delayed_u0=1'h0;
reg	[15:0]	syncEnable_u29=16'h0;
reg		reg_644a10e2_result_delayed_result_delayed_u0=1'h0;
reg	[15:0]	syncEnable_u30_u0=16'h0;
assign simplePinWrite=GO&{1{GO}};
assign and_u641_u0=done_cache_u40&port_0ba14e5d_;
assign or_u168_u0=and_u641_u0|RESET;
always @(posedge CLK or posedge GO or posedge or_u168_u0)
begin
if (or_u168_u0)
done_cache_u40<=1'h0;
else if (GO)
done_cache_u40<=1'h1;
else done_cache_u40<=done_cache_u40;
end
assign and_u646_u0=done_cache_u41_u0&port_0ba14e5d_;
always @(posedge CLK or posedge reg_644a10e2_u0 or posedge or_u169_u0)
begin
if (or_u169_u0)
done_cache_u41_u0<=1'h0;
else if (reg_644a10e2_u0)
done_cache_u41_u0<=1'h1;
else done_cache_u41_u0<=done_cache_u41_u0;
end
assign or_u169_u0=and_u646_u0|RESET;
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_7779df0d_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_7779df0d_instance(.GO(reg_644a10e2_result_delayed_u0), 
  .port_661c2da4_(syncEnable_u29), .port_0186947a_(port_610b7aeb_), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_7779df0d_instance_RESULT));
always @(posedge CLK or posedge reg_6857eec0_u0 or posedge or_u170_u0)
begin
if (or_u170_u0)
reg_663425d2_u0<=1'h0;
else if (reg_6857eec0_u0)
reg_663425d2_u0<=1'h1;
else reg_663425d2_u0<=reg_663425d2_u0;
end
assign and_u655_u0=reg_663425d2_u0&port_0ba14e5d_;
assign or_u170_u0=and_u655_u0|RESET;
assign add=port_5330dddc_+32'h1;
assign add_u11=port_0e198730_+16'h1;
assign not_u125=!port_55a91fbd_;
assign simplePinWrite_u102=reg_644a10e2_result_delayed_u0&{1{reg_644a10e2_result_delayed_u0}};
assign simplePinWrite_u103=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_7779df0d_instance_RESULT&{16{reg_644a10e2_result_delayed_u0}};
assign simplePinWrite_u104=16'h1&{16{1'h1}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7fa5a9ca_u0<=1'h0;
else reg_7fa5a9ca_u0<=reg_6857eec0_u0;
end
assign or_u171_u0=GO|reg_644a10e2_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6857eec0_u0<=1'h0;
else reg_6857eec0_u0<=reg_644a10e2_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_644a10e2_u0<=1'h0;
else reg_644a10e2_u0<=reg_5a7b2b71_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5a7b2b71_u0<=1'h0;
else reg_5a7b2b71_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_644a10e2_result_delayed_u0<=1'h0;
else reg_644a10e2_result_delayed_u0<=reg_644a10e2_u0;
end
always @(posedge CLK)
begin
if (reg_5a7b2b71_u0)
syncEnable_u29<=port_610b7aeb_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_644a10e2_result_delayed_result_delayed_u0<=1'h0;
else reg_644a10e2_result_delayed_result_delayed_u0<=reg_644a10e2_result_delayed_u0;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u30_u0<=port_58e85b4e_;
end
assign RESULT=GO;
assign RESULT_u355=16'h0;
assign RESULT_u356=GO;
assign RESULT_u357=add;
assign RESULT_u358=GO;
assign RESULT_u359=add_u11;
assign RESULT_u360=GO;
assign RESULT_u361=16'h0;
assign RESULT_u362=GO;
assign RESULT_u363=not_u125;
assign RESULT_u364=or_u171_u0;
assign RESULT_u365=32'h0;
assign RESULT_u366=3'h1;
assign RESULT_u367=reg_6857eec0_u0;
assign RESULT_u368=32'h0;
assign RESULT_u369=syncEnable_u30_u0;
assign RESULT_u370=3'h1;
assign RESULT_u371=simplePinWrite;
assign RESULT_u372=simplePinWrite_u104;
assign RESULT_u373=simplePinWrite_u102;
assign RESULT_u374=simplePinWrite_u103;
assign DONE=reg_7fa5a9ca_u0;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_7779df0d_(GO, port_661c2da4_, port_0186947a_, RESULT);
input		GO;
input	[15:0]	port_661c2da4_;
input	[15:0]	port_0186947a_;
output	[15:0]	RESULT;
wire	[16:0]	add;
wire	[15:0]	LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_2fb496b7_instance_RESULT;
assign add={port_661c2da4_[15], port_661c2da4_}+{port_0186947a_[15], port_0186947a_};
LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_2fb496b7_ LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_2fb496b7_instance(.GO(GO), 
  .port_6db40575_({add[16], add[16:2]}), .RESULT(LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_2fb496b7_instance_RESULT));
assign RESULT=LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_2fb496b7_instance_RESULT;
endmodule



module LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_LL1_H_iunzipFilter2D_procedure_2fb496b7_(GO, port_6db40575_, RESULT);
input		GO;
input	[15:0]	port_6db40575_;
output	[15:0]	RESULT;
wire		greaterThan;
wire signed	[15:0]	greaterThan_a_signed;
wire signed	[15:0]	greaterThan_b_signed;
wire		not_u124_u0;
wire		and_u650_u0;
wire		and_u651_u0;
wire		and_u652_u0;
wire	[15:0]	mux_u43;
wire		and_u653_u0;
assign greaterThan_a_signed=16'h0;
assign greaterThan_b_signed=port_6db40575_;
assign greaterThan=greaterThan_a_signed>greaterThan_b_signed;
assign not_u124_u0=~greaterThan;
assign and_u650_u0=GO&not_u124_u0;
assign and_u651_u0=GO&greaterThan;
assign and_u652_u0=and_u651_u0&GO;
assign mux_u43=(and_u652_u0)?16'h0:port_6db40575_;
assign and_u653_u0=and_u650_u0&GO;
assign RESULT=mux_u43;
endmodule


