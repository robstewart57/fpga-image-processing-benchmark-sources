// __  ___ __ ___  _ __   ___  ___ 
// \ \/ / '__/ _ \| '_ \ / _ \/ __|
//  >  <| | | (_) | | | | (_) \__ \
// /_/\_\_|  \___/|_| |_|\___/|___/
// 
// Xronos synthesizer version
// Run date: Thu 2 Nov 2017 13:59:44 +0000
// 

module resized_LH3_xy(Out1_SEND, Out1_ACK, Out1_DATA, Out1_RDY, Out1_COUNT, In1_ACK, In1_COUNT, RESET, CLK, In1_SEND, In1_DATA);
output		Out1_SEND;
input		Out1_ACK;
wire		consumeRow_done;
wire		reset_done;
wire		repeatRowExpanded_go;
output	[15:0]	Out1_DATA;
input		Out1_RDY;
wire		reset_go;
output	[15:0]	Out1_COUNT;
output		In1_ACK;
input	[15:0]	In1_COUNT;
input		RESET;
wire		repeatRowExpanded_done;
input		CLK;
input		In1_SEND;
wire		consumeRow_go;
input	[15:0]	In1_DATA;
wire	[15:0]	scheduler_u344;
wire	[15:0]	scheduler_u346;
wire		scheduler_u348;
wire	[31:0]	scheduler_u338;
wire		resized_LH3_xy_scheduler_instance_DONE;
wire	[31:0]	scheduler_u332;
wire		scheduler_u345;
wire	[2:0]	scheduler_u343;
wire		scheduler_u333;
wire		scheduler_u337;
wire		scheduler_u340;
wire	[31:0]	scheduler_u336;
wire		scheduler_u334;
wire		scheduler_u349;
wire	[31:0]	scheduler_u342;
wire		scheduler;
wire		scheduler_u339;
wire		scheduler_u347;
wire		scheduler_u335;
wire		scheduler_u341;
wire		bus_01b00d94_;
wire		bus_5cd62f8e_;
wire	[15:0]	bus_6f4f27ab_;
wire	[15:0]	bus_0859aa58_;
wire	[31:0]	bus_1598a4d3_;
wire		bus_4eb99653_;
wire		bus_39892bbf_;
wire	[15:0]	bus_7927363a_;
wire	[2:0]	bus_1310b3e4_;
wire		bus_604acdab_;
wire		bus_4497015b_;
wire		bus_5d365df5_;
wire		bus_45a18503_;
wire		bus_3606f0fa_;
wire		bus_7223468d_;
wire	[15:0]	bus_33af6980_;
wire	[15:0]	bus_5e36be26_;
wire		bus_3866f699_;
wire	[31:0]	bus_48c16de3_;
wire	[31:0]	bus_36c9b0d0_;
wire		bus_38031f96_;
wire	[15:0]	bus_07b29725_;
wire	[15:0]	bus_21d6a5fd_;
wire		bus_30f6e3b0_;
wire		bus_12a86ec5_;
wire	[2:0]	bus_6620e554_;
wire		bus_2f725b02_;
wire		bus_61fe06bb_;
wire		repeatRowExpanded;
wire		repeatRowExpanded_u44;
wire	[15:0]	repeatRowExpanded_u46;
wire	[2:0]	repeatRowExpanded_u43;
wire		resized_LH3_xy_repeatRowExpanded_instance_DONE;
wire	[31:0]	repeatRowExpanded_u42;
wire	[31:0]	repeatRowExpanded_u45;
wire	[15:0]	repeatRowExpanded_u40;
wire		repeatRowExpanded_u41;
wire	[2:0]	repeatRowExpanded_u47;
wire	[31:0]	bus_32281ea7_;
wire		reset_u16;
wire		resized_LH3_xy_reset_instance_DONE;
wire	[15:0]	reset_u17;
wire		reset;
wire	[15:0]	reset_u15;
wire	[31:0]	bus_14dbd04d_;
wire		bus_07319e33_;
wire	[2:0]	consumeRow_u54;
wire	[31:0]	consumeRow_u52;
wire	[15:0]	consumeRow_u53;
wire	[2:0]	consumeRow_u58;
wire	[15:0]	consumeRow_u57;
wire	[15:0]	consumeRow_u50;
wire		consumeRow_u59;
wire	[31:0]	consumeRow_u56;
wire		consumeRow;
wire		resized_LH3_xy_consumeRow_instance_DONE;
wire		consumeRow_u51;
wire		consumeRow_u55;
wire		bus_2186a09b_;
wire	[15:0]	bus_04fa5f53_;
assign Out1_SEND=scheduler_u345;
assign consumeRow_done=bus_01b00d94_;
assign reset_done=bus_3866f699_;
assign repeatRowExpanded_go=scheduler_u348;
assign Out1_DATA=scheduler_u346;
assign reset_go=scheduler_u349;
assign Out1_COUNT=scheduler_u344;
assign In1_ACK=consumeRow_u59;
assign repeatRowExpanded_done=bus_7223468d_;
assign consumeRow_go=scheduler_u347;
resized_LH3_xy_scheduler resized_LH3_xy_scheduler_instance(.CLK(CLK), .RESET(bus_45a18503_), 
  .GO(bus_3606f0fa_), .port_3a102d1f_(32'h0), .port_6cb7d4b7_(bus_61fe06bb_), .port_639e94f2_(bus_32281ea7_), 
  .port_072ed7ee_(bus_14dbd04d_), .port_202620a3_(bus_07319e33_), .port_1bba0a1c_(bus_33af6980_), 
  .port_4c65738f_(bus_5e36be26_), .port_03915889_(bus_4eb99653_), .port_5c53ee9c_(bus_0859aa58_), 
  .port_7fb2b3af_(Out1_RDY), .port_4f7d225f_(repeatRowExpanded_done), .port_157e6b5b_(In1_SEND), 
  .port_13873765_(consumeRow_done), .port_56dbc9e6_(reset_done), .DONE(resized_LH3_xy_scheduler_instance_DONE), 
  .RESULT(scheduler), .RESULT_u2370(scheduler_u332), .RESULT_u2371(scheduler_u333), 
  .RESULT_u2372(scheduler_u334), .RESULT_u2373(scheduler_u335), .RESULT_u2374(scheduler_u336), 
  .RESULT_u2375(scheduler_u337), .RESULT_u2376(scheduler_u338), .RESULT_u2377(scheduler_u339), 
  .RESULT_u2378(scheduler_u340), .RESULT_u2379(scheduler_u341), .RESULT_u2380(scheduler_u342), 
  .RESULT_u2381(scheduler_u343), .RESULT_u2382(scheduler_u344), .RESULT_u2383(scheduler_u345), 
  .RESULT_u2384(scheduler_u346), .RESULT_u2385(scheduler_u347), .RESULT_u2386(scheduler_u348), 
  .RESULT_u2387(scheduler_u349));
assign bus_01b00d94_=resized_LH3_xy_consumeRow_instance_DONE&{1{resized_LH3_xy_consumeRow_instance_DONE}};
resized_LH3_xy_structuralmemory_5a4854c1_ resized_LH3_xy_structuralmemory_5a4854c1__1(.CLK_u23(CLK), 
  .bus_4424cad2_(bus_45a18503_), .bus_287c41c7_(bus_36c9b0d0_), .bus_66538fba_(3'h1), 
  .bus_793de9c2_(bus_30f6e3b0_), .bus_1f47f383_(bus_2f725b02_), .bus_462ad95f_(bus_07b29725_), 
  .bus_6f4f27ab_(bus_6f4f27ab_), .bus_5cd62f8e_(bus_5cd62f8e_));
resized_LH3_xy_simplememoryreferee_4dbf2a2f_ resized_LH3_xy_simplememoryreferee_4dbf2a2f__1(.bus_170ffe51_(CLK), 
  .bus_2bdc80e5_(bus_45a18503_), .bus_5068a6cf_(bus_2186a09b_), .bus_4a24c1e1_(bus_04fa5f53_), 
  .bus_71489945_(consumeRow_u55), .bus_0668b190_(consumeRow_u57), .bus_69dc047c_(consumeRow_u56), 
  .bus_419996e9_(3'h1), .bus_309461d8_(repeatRowExpanded_u44), .bus_0943531d_(repeatRowExpanded_u46), 
  .bus_1bce23d3_(repeatRowExpanded_u45), .bus_6d8c43ff_(3'h1), .bus_67ef8aa5_(scheduler_u341), 
  .bus_3032e61d_(scheduler_u342), .bus_7a45fad8_(3'h1), .bus_7927363a_(bus_7927363a_), 
  .bus_1598a4d3_(bus_1598a4d3_), .bus_39892bbf_(bus_39892bbf_), .bus_604acdab_(bus_604acdab_), 
  .bus_1310b3e4_(bus_1310b3e4_), .bus_4497015b_(bus_4497015b_), .bus_5d365df5_(bus_5d365df5_), 
  .bus_0859aa58_(bus_0859aa58_), .bus_4eb99653_(bus_4eb99653_));
resized_LH3_xy_globalreset_physical_6b469655_ resized_LH3_xy_globalreset_physical_6b469655__1(.bus_7bfcb29f_(CLK), 
  .bus_21c9004a_(RESET), .bus_45a18503_(bus_45a18503_));
resized_LH3_xy_Kicker_47 resized_LH3_xy_Kicker_47_1(.CLK(CLK), .RESET(bus_45a18503_), 
  .bus_3606f0fa_(bus_3606f0fa_));
assign bus_7223468d_=resized_LH3_xy_repeatRowExpanded_instance_DONE&{1{resized_LH3_xy_repeatRowExpanded_instance_DONE}};
resized_LH3_xy_stateVar_x resized_LH3_xy_stateVar_x_1(.bus_21f26c1b_(CLK), .bus_27078042_(bus_45a18503_), 
  .bus_318dd820_(consumeRow), .bus_18336d09_(consumeRow_u50), .bus_26bd9abe_(reset_u16), 
  .bus_49e109b4_(16'h0), .bus_33af6980_(bus_33af6980_));
resized_LH3_xy_stateVar_rowRepeated resized_LH3_xy_stateVar_rowRepeated_1(.bus_45f031f5_(CLK), 
  .bus_1b617bad_(bus_45a18503_), .bus_3bba85fa_(repeatRowExpanded), .bus_6fadc4af_(repeatRowExpanded_u40), 
  .bus_4ba53be4_(reset), .bus_3e7ecbe0_(16'h1), .bus_5e36be26_(bus_5e36be26_));
assign bus_3866f699_=resized_LH3_xy_reset_instance_DONE&{1{resized_LH3_xy_reset_instance_DONE}};
resized_LH3_xy_stateVar_fsmOldState_resized_LH3_xy resized_LH3_xy_stateVar_fsmOldState_resized_LH3_xy_1(.bus_1e850958_(CLK), 
  .bus_0fe2bf8a_(bus_45a18503_), .bus_2d9446c1_(scheduler), .bus_0169b7ea_(32'h0), 
  .bus_48c16de3_(bus_48c16de3_));
resized_LH3_xy_simplememoryreferee_10f2e65e_ resized_LH3_xy_simplememoryreferee_10f2e65e__1(.bus_095cf1de_(CLK), 
  .bus_1d16e5f4_(bus_45a18503_), .bus_15440525_(bus_5cd62f8e_), .bus_1f52af7b_(bus_6f4f27ab_), 
  .bus_5d57546f_(consumeRow_u51), .bus_23881311_(consumeRow_u53), .bus_385fd4fe_(consumeRow_u52), 
  .bus_074a4e9c_(3'h1), .bus_0109f5e5_(repeatRowExpanded_u41), .bus_38ee4680_(repeatRowExpanded_u42), 
  .bus_55728af0_(3'h1), .bus_07b29725_(bus_07b29725_), .bus_36c9b0d0_(bus_36c9b0d0_), 
  .bus_2f725b02_(bus_2f725b02_), .bus_30f6e3b0_(bus_30f6e3b0_), .bus_6620e554_(bus_6620e554_), 
  .bus_38031f96_(bus_38031f96_), .bus_21d6a5fd_(bus_21d6a5fd_), .bus_12a86ec5_(bus_12a86ec5_));
resized_LH3_xy_stateVar_fsmState_resized_LH3_xy resized_LH3_xy_stateVar_fsmState_resized_LH3_xy_1(.bus_35a4b222_(CLK), 
  .bus_1fa30b0d_(bus_45a18503_), .bus_7894e09d_(scheduler_u333), .bus_6f4dfd67_(scheduler_u334), 
  .bus_61fe06bb_(bus_61fe06bb_));
resized_LH3_xy_repeatRowExpanded resized_LH3_xy_repeatRowExpanded_instance(.CLK(CLK), 
  .RESET(bus_45a18503_), .GO(repeatRowExpanded_go), .port_7ef0238d_(bus_5e36be26_), 
  .port_183b6d71_(bus_12a86ec5_), .port_466e1c3e_(bus_21d6a5fd_), .port_138273d0_(bus_5d365df5_), 
  .DONE(resized_LH3_xy_repeatRowExpanded_instance_DONE), .RESULT(repeatRowExpanded), 
  .RESULT_u2388(repeatRowExpanded_u40), .RESULT_u2393(repeatRowExpanded_u41), 
  .RESULT_u2394(repeatRowExpanded_u42), .RESULT_u2395(repeatRowExpanded_u43), 
  .RESULT_u2389(repeatRowExpanded_u44), .RESULT_u2390(repeatRowExpanded_u45), 
  .RESULT_u2391(repeatRowExpanded_u46), .RESULT_u2392(repeatRowExpanded_u47));
resized_LH3_xy_stateVar_Out1TokenIndex resized_LH3_xy_stateVar_Out1TokenIndex_1(.bus_240b7571_(CLK), 
  .bus_2effa3d4_(bus_45a18503_), .bus_69e423e6_(scheduler_u335), .bus_45898356_(scheduler_u336), 
  .bus_32281ea7_(bus_32281ea7_));
resized_LH3_xy_reset resized_LH3_xy_reset_instance(.CLK(CLK), .RESET(bus_45a18503_), 
  .GO(reset_go), .DONE(resized_LH3_xy_reset_instance_DONE), .RESULT(reset), .RESULT_u2396(reset_u15), 
  .RESULT_u2397(reset_u16), .RESULT_u2398(reset_u17));
resized_LH3_xy_stateVar_Out1MaxTokenIndex resized_LH3_xy_stateVar_Out1MaxTokenIndex_1(.bus_7dd8451b_(CLK), 
  .bus_6e8b3703_(bus_45a18503_), .bus_185d6703_(scheduler_u337), .bus_10961150_(scheduler_u338), 
  .bus_14dbd04d_(bus_14dbd04d_));
resized_LH3_xy_stateVar_Out1PortEnable resized_LH3_xy_stateVar_Out1PortEnable_1(.bus_66c9187f_(CLK), 
  .bus_7bb89c8a_(bus_45a18503_), .bus_016a15f2_(scheduler_u339), .bus_10ad7aff_(scheduler_u340), 
  .bus_07319e33_(bus_07319e33_));
resized_LH3_xy_consumeRow resized_LH3_xy_consumeRow_instance(.CLK(CLK), .RESET(bus_45a18503_), 
  .GO(consumeRow_go), .port_7ee25a17_(bus_33af6980_), .port_4bf12c4e_(bus_38031f96_), 
  .port_00eaa84f_(bus_4497015b_), .port_0266fa2c_(In1_DATA), .DONE(resized_LH3_xy_consumeRow_instance_DONE), 
  .RESULT(consumeRow), .RESULT_u2399(consumeRow_u50), .RESULT_u2404(consumeRow_u51), 
  .RESULT_u2405(consumeRow_u52), .RESULT_u2406(consumeRow_u53), .RESULT_u2407(consumeRow_u54), 
  .RESULT_u2400(consumeRow_u55), .RESULT_u2401(consumeRow_u56), .RESULT_u2402(consumeRow_u57), 
  .RESULT_u2403(consumeRow_u58), .RESULT_u2408(consumeRow_u59));
resized_LH3_xy_structuralmemory_46badd45_ resized_LH3_xy_structuralmemory_46badd45__1(.CLK_u24(CLK), 
  .bus_568ab95c_(bus_45a18503_), .bus_12817703_(bus_1598a4d3_), .bus_12f2a754_(3'h1), 
  .bus_1cfe3bb9_(bus_604acdab_), .bus_183866fe_(bus_39892bbf_), .bus_6170e247_(bus_7927363a_), 
  .bus_04fa5f53_(bus_04fa5f53_), .bus_2186a09b_(bus_2186a09b_));
endmodule



module resized_LH3_xy_scheduler(CLK, RESET, GO, port_3a102d1f_, port_6cb7d4b7_, port_639e94f2_, port_072ed7ee_, port_202620a3_, port_1bba0a1c_, port_4c65738f_, port_03915889_, port_5c53ee9c_, port_7fb2b3af_, port_4f7d225f_, port_157e6b5b_, port_13873765_, port_56dbc9e6_, RESULT, RESULT_u2370, RESULT_u2371, RESULT_u2372, RESULT_u2373, RESULT_u2374, RESULT_u2375, RESULT_u2376, RESULT_u2377, RESULT_u2378, RESULT_u2379, RESULT_u2380, RESULT_u2381, RESULT_u2382, RESULT_u2383, RESULT_u2384, RESULT_u2385, RESULT_u2386, RESULT_u2387, DONE);
input		CLK;
input		RESET;
input		GO;
input	[31:0]	port_3a102d1f_;
input		port_6cb7d4b7_;
input	[31:0]	port_639e94f2_;
input	[31:0]	port_072ed7ee_;
input		port_202620a3_;
input	[15:0]	port_1bba0a1c_;
input	[15:0]	port_4c65738f_;
input		port_03915889_;
input	[15:0]	port_5c53ee9c_;
input		port_7fb2b3af_;
input		port_4f7d225f_;
input		port_157e6b5b_;
input		port_13873765_;
input		port_56dbc9e6_;
output		RESULT;
output	[31:0]	RESULT_u2370;
output		RESULT_u2371;
output		RESULT_u2372;
output		RESULT_u2373;
output	[31:0]	RESULT_u2374;
output		RESULT_u2375;
output	[31:0]	RESULT_u2376;
output		RESULT_u2377;
output		RESULT_u2378;
output		RESULT_u2379;
output	[31:0]	RESULT_u2380;
output	[2:0]	RESULT_u2381;
output	[15:0]	RESULT_u2382;
output		RESULT_u2383;
output	[15:0]	RESULT_u2384;
output		RESULT_u2385;
output		RESULT_u2386;
output		RESULT_u2387;
output		DONE;
wire	[15:0]	lessThan_b_unsigned;
wire		lessThan;
wire	[15:0]	lessThan_a_unsigned;
wire		equals;
wire	[15:0]	equals_a_unsigned;
wire	[15:0]	equals_b_unsigned;
wire	[15:0]	lessThan_u98_b_unsigned;
wire	[15:0]	lessThan_u98_a_unsigned;
wire		lessThan_u98;
wire		andOp;
wire	[15:0]	equals_u212_a_unsigned;
wire		equals_u212;
wire	[15:0]	equals_u212_b_unsigned;
wire signed	[31:0]	equals_u213_a_signed;
wire		equals_u213;
wire signed	[31:0]	equals_u213_b_signed;
wire		not_u645_u0;
wire		and_u4058_u0;
wire		and_u4059_u0;
wire		andOp_u213;
wire		and_u4060_u0;
wire		not_u646_u0;
wire		and_u4061_u0;
wire		simplePinWrite;
wire		not_u647_u0;
wire		and_u4062_u0;
wire		and_u4063_u0;
wire		simplePinWrite_u566;
wire		and_u4064_u0;
wire		not_u648_u0;
wire		and_u4065_u0;
wire		simplePinWrite_u567;
wire		and_u4066_u0;
reg		reg_4985bd85_u0=1'h0;
reg		reg_35c809c8_u0=1'h0;
reg		reg_5760cf63_u0=1'h0;
reg		reg_6fb08fb4_u0=1'h0;
reg		reg_4ff7f3f0_u0=1'h0;
reg		reg_3027d020_u0=1'h0;
reg		reg_794edd46_u0=1'h0;
reg		reg_3726932e_u0=1'h0;
reg		reg_3d184510_u0=1'h0;
reg		reg_59d7b5da_u0=1'h0;
reg		reg_16604e6f_u0=1'h0;
reg		reg_6903fd17_u0=1'h0;
reg		reg_7aa64abe_u0=1'h0;
reg		reg_1885f09c_u0=1'h0;
reg		reg_2faca78c_u0=1'h0;
reg		reg_57323713_u0=1'h0;
reg		reg_20d1a0f8_u0=1'h0;
reg		reg_20d7d0fd_u0=1'h0;
reg		reg_4787c3ad_u0=1'h0;
reg		reg_4274ae45_u0=1'h0;
reg		reg_2b115723_u0=1'h0;
reg		reg_330dd339_u0=1'h0;
reg		reg_6aa30297_u0=1'h0;
reg		reg_45ddb9e8_u0=1'h0;
reg		reg_594f457a_u0=1'h0;
reg		reg_74b6d880_u0=1'h0;
reg		reg_4490a0a8_u0=1'h0;
reg		reg_3cb65c8f_u0=1'h0;
reg		reg_0dbaa983_u0=1'h0;
reg		reg_45c4b9fe_u0=1'h0;
reg		reg_21729149_u0=1'h0;
reg		reg_3c7ba446_u0=1'h0;
reg		reg_1b5e971f_u0=1'h0;
reg		reg_36d13294_u0=1'h0;
reg		reg_210fdd48_u0=1'h0;
reg		reg_45e011aa_u0=1'h0;
reg		reg_21729149_result_delayed_u0=1'h0;
reg		reg_55e64da9_u0=1'h0;
reg		reg_19fcf5ae_u0=1'h0;
reg		reg_0858480b_u0=1'h0;
reg		reg_21729149_result_delayed_result_delayed_u0=1'h0;
reg		reg_6ceba0be_u0=1'h0;
reg		reg_068d86d5_u0=1'h0;
reg		reg_746c5835_u0=1'h0;
reg		reg_0672d22b_u0=1'h0;
reg		reg_3d3b0167_u0=1'h0;
reg		reg_55e64da9_result_delayed_u0=1'h0;
reg		reg_343be065_u0=1'h0;
reg		reg_145a1005_u0=1'h0;
reg		reg_4cbad8e5_u0=1'h0;
reg		reg_42c646a7_u0=1'h0;
reg		reg_5e145a76_u0=1'h0;
reg		reg_63b54bd2_u0=1'h0;
reg		reg_29b64ddf_u0=1'h0;
reg		reg_0120594a_u0=1'h0;
reg		reg_049c34f3_u0=1'h0;
reg		reg_244f643a_u0=1'h0;
reg		reg_49a5b9d0_u0=1'h0;
reg		reg_741cf86b_u0=1'h0;
reg		reg_0e961ae8_u0=1'h0;
reg		reg_728c76f2_u0=1'h0;
reg		reg_0e961ae8_result_delayed_u0=1'h0;
reg		reg_37142796_u0=1'h0;
reg		reg_4cae982d_u0=1'h0;
reg		reg_6b924716_u0=1'h0;
reg		reg_7ad2c256_u0=1'h0;
reg		reg_413e1dbb_u0=1'h0;
reg		reg_3f89f30c_u0=1'h0;
reg		reg_44c1644a_u0=1'h0;
reg		reg_3e622eee_u0=1'h0;
reg		reg_39988114_u0=1'h0;
reg		reg_16a5622b_u0=1'h0;
reg		reg_5f70cbfe_u0=1'h0;
reg		reg_7a53eec3_u0=1'h0;
reg		reg_2d178d82_u0=1'h0;
reg		reg_50958802_u0=1'h0;
reg		reg_430f0398_u0=1'h0;
reg		reg_67e7177f_u0=1'h0;
reg		reg_06c0f659_u0=1'h0;
reg		reg_210fdd48_result_delayed_u0=1'h0;
reg		reg_14042498_u0=1'h0;
reg		reg_6b03bf9f_u0=1'h0;
reg		reg_7e53b6cf_u0=1'h0;
reg		reg_0d002d9e_u0=1'h0;
reg		reg_2927f9b8_u0=1'h0;
reg		reg_4dc3c160_u0=1'h0;
reg		reg_37a25b06_u0=1'h0;
reg		reg_473d6b97_u0=1'h0;
reg		reg_068d86d5_result_delayed_u0=1'h0;
reg		reg_550541a9_u0=1'h0;
reg		reg_3131c19c_u0=1'h0;
reg		reg_6f4947f8_u0=1'h0;
reg		reg_16604e6f_result_delayed_u0=1'h0;
reg		reg_2b76cbc2_u0=1'h0;
reg		reg_09925d27_u0=1'h0;
reg		reg_00ca0473_u0=1'h0;
reg		reg_63b54bd2_result_delayed_u0=1'h0;
reg		reg_69c13d7a_u0=1'h0;
reg		reg_5f70cbfe_result_delayed_u0=1'h0;
reg		reg_14ea9829_u0=1'h0;
reg		reg_24743cb0_u0=1'h0;
reg		reg_75f8153e_u0=1'h0;
reg		reg_6b924716_result_delayed_u0=1'h0;
reg		reg_2339dbf0_u0=1'h0;
reg		reg_11bc6171_u0=1'h0;
reg		reg_6af44a24_u0=1'h0;
reg		reg_0c1a90ca_u0=1'h0;
reg		reg_4a3d5eec_u0=1'h0;
reg		reg_2339dbf0_result_delayed_u0=1'h0;
reg		reg_29b64ddf_result_delayed_u0=1'h0;
reg		reg_0858480b_result_delayed_u0=1'h0;
reg		reg_2eca9a1d_u0=1'h0;
reg		reg_142e74f6_u0=1'h0;
reg		reg_7bcb7712_u0=1'h0;
reg		reg_37f5df2f_u0=1'h0;
reg		reg_2b76cbc2_result_delayed_u0=1'h0;
reg		reg_6da5dd78_u0=1'h0;
reg		reg_794edd46_result_delayed_u0=1'h0;
reg		reg_29875567_u0=1'h0;
reg		reg_55e64da9_result_delayed_result_delayed_u0=1'h0;
reg		reg_393565d7_u0=1'h0;
reg		reg_3b51abb4_u0=1'h0;
reg		reg_21f11516_u0=1'h0;
reg		reg_41b4a953_u0=1'h0;
reg		reg_671babf3_u0=1'h0;
reg		reg_3a57c6ba_u0=1'h0;
reg		reg_6afd820d_u0=1'h0;
reg		reg_393565d7_result_delayed_u0=1'h0;
reg		reg_6d8fa179_u0=1'h0;
reg		reg_19be9d49_u0=1'h0;
reg		reg_7a61a699_u0=1'h0;
reg		reg_1dad4554_u0=1'h0;
reg		reg_3a5d4aa0_u0=1'h0;
reg		reg_660f9ef1_u0=1'h0;
reg		reg_1f3d8a38_u0=1'h0;
reg		reg_430f0398_result_delayed_u0=1'h0;
reg		reg_7aa64abe_result_delayed_u0=1'h0;
reg		reg_210fdd48_result_delayed_result_delayed_u0=1'h0;
reg		reg_2e9f4b96_u0=1'h0;
reg		reg_7d2bf821_u0=1'h0;
reg		reg_5760cf63_result_delayed_u0=1'h0;
reg		reg_2eca9a1d_result_delayed_u0=1'h0;
reg		reg_3c50cd45_u0=1'h0;
reg		reg_4cae982d_result_delayed_u0=1'h0;
reg		reg_07c27ed5_u0=1'h0;
reg		reg_1f3d8a38_result_delayed_u0=1'h0;
reg		reg_1a329b29_u0=1'h0;
reg		reg_4d3f2823_u0=1'h0;
reg		reg_4f36662b_u0=1'h0;
reg		reg_3fe03efe_u0=1'h0;
reg		reg_75f2c8ed_u0=1'h0;
reg		reg_3c0ef12e_u0=1'h0;
reg		reg_3c568577_u0=1'h0;
reg		reg_1885f09c_result_delayed_u0=1'h0;
reg		reg_2c201504_u0=1'h0;
reg		reg_618a90a2_u0=1'h0;
reg		reg_5e145a76_result_delayed_u0=1'h0;
reg		reg_618a90a2_result_delayed_u0=1'h0;
reg		reg_64d83df2_u0=1'h0;
reg		reg_594f457a_result_delayed_u0=1'h0;
reg		reg_7aa64abe_result_delayed_result_delayed_u0=1'h0;
reg		reg_529137a1_u0=1'h0;
reg		reg_53e492d4_u0=1'h0;
reg		reg_0833f502_u0=1'h0;
reg		reg_1b5e971f_result_delayed_u0=1'h0;
reg		reg_0c1a90ca_result_delayed_u0=1'h0;
reg		reg_142e74f6_result_delayed_u0=1'h0;
reg		reg_07f782c9_u0=1'h0;
reg		reg_1980ccbe_u0=1'h0;
reg		reg_63b54bd2_result_delayed_result_delayed_u0=1'h0;
reg		reg_45c4b9fe_result_delayed_u0=1'h0;
reg		reg_3d3b0167_result_delayed_u0=1'h0;
reg		reg_6af44a24_result_delayed_u0=1'h0;
reg		reg_6abcb3ff_u0=1'h0;
reg		reg_6d25a062_u0=1'h0;
reg		reg_48d7a190_u0=1'h0;
wire		mux_u404;
wire		or_u1205_u0;
reg		reg_4b73b23b_u0=1'h0;
reg		reg_22e61fae_u0=1'h0;
reg		reg_69dda494_u0=1'h0;
reg		reg_3cbd59f7_u0=1'h0;
reg		reg_0e9d33d1_u0=1'h0;
reg		reg_2d8038cc_u0=1'h0;
reg		reg_7213e342_u0=1'h0;
reg		reg_222a4f78_u0=1'h0;
reg		reg_0dbaa983_result_delayed_u0=1'h0;
reg		reg_3c50cd45_result_delayed_u0=1'h0;
reg		reg_56f347a4_u0=1'h0;
reg		reg_01dd2487_u0=1'h0;
reg		reg_238aead6_u0=1'h0;
reg		reg_5a3ed760_u0=1'h0;
reg		reg_79d4808b_u0=1'h0;
reg		reg_6fb08fb4_result_delayed_u0=1'h0;
reg		reg_3d184510_result_delayed_u0=1'h0;
reg		reg_430f0398_result_delayed_result_delayed_u0=1'h0;
reg		reg_6535b053_u0=1'h0;
reg		reg_7aa64abe_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_6d25a062_result_delayed_u0=1'h0;
reg		reg_618a90a2_result_delayed_result_delayed_u0=1'h0;
reg		reg_79c318b3_u0=1'h0;
reg		reg_28ebf99a_u0=1'h0;
reg		reg_2376da04_u0=1'h0;
reg		reg_512aac58_u0=1'h0;
reg		reg_5091b5e2_u0=1'h0;
reg		reg_741cf86b_result_delayed_u0=1'h0;
reg		reg_6abcb3ff_result_delayed_u0=1'h0;
reg		reg_46861ff1_u0=1'h0;
reg		reg_3131c19c_result_delayed_u0=1'h0;
reg		reg_0269f3e8_u0=1'h0;
reg		reg_1b5e971f_result_delayed_result_delayed_u0=1'h0;
reg		reg_23129694_u0=1'h0;
reg		reg_6aa9532f_u0=1'h0;
reg		reg_2a0b1f83_u0=1'h0;
reg		reg_07b96631_u0=1'h0;
reg		reg_517738fd_u0=1'h0;
reg		reg_42c646a7_result_delayed_u0=1'h0;
reg		reg_01dd2487_result_delayed_u0=1'h0;
reg		reg_242dc5a0_u0=1'h0;
reg		reg_003f51b2_u0=1'h0;
reg		reg_2cb66d26_u0=1'h0;
reg		reg_794edd46_result_delayed_result_delayed_u0=1'h0;
reg		reg_309c310d_u0=1'h0;
reg		reg_0a6b2ffa_u0=1'h0;
wire		and_u4067_u0;
reg		reg_517738fd_result_delayed_u0=1'h0;
reg		reg_358f4c1c_u0=1'h0;
reg		reg_7ad08748_u0=1'h0;
reg		reg_320deb94_u0=1'h0;
reg		reg_60829d18_u0=1'h0;
reg		reg_395b58c5_u0=1'h0;
reg		reg_222c2bb3_u0=1'h0;
reg		reg_57323713_result_delayed_u0=1'h0;
reg		reg_7101c0a1_u0=1'h0;
reg		reg_550d08a9_u0=1'h0;
reg		reg_6903fd17_result_delayed_u0=1'h0;
reg		reg_2faca78c_result_delayed_u0=1'h0;
reg		reg_343be065_result_delayed_u0=1'h0;
reg		reg_73be9a15_u0=1'h0;
reg		reg_7213e342_result_delayed_u0=1'h0;
reg		reg_2f1102bc_u0=1'h0;
reg		reg_3cb65c8f_result_delayed_u0=1'h0;
reg		reg_7aa64abe_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_4977a8c0_u0=1'h0;
reg		reg_2c201504_result_delayed_u0=1'h0;
reg		reg_4cbad8e5_result_delayed_u0=1'h0;
reg		reg_06c0f659_result_delayed_u0=1'h0;
reg		reg_6d8fa179_result_delayed_u0=1'h0;
reg		reg_29875567_result_delayed_u0=1'h0;
reg		reg_4beb2654_u0=1'h0;
reg		reg_4ee47324_u0=1'h0;
reg		reg_3a3faffe_u0=1'h0;
reg		reg_79d4808b_result_delayed_u0=1'h0;
reg		reg_24743cb0_result_delayed_u0=1'h0;
reg		reg_343be065_result_delayed_result_delayed_u0=1'h0;
reg		reg_5ec29f05_u0=1'h0;
reg		reg_4985bd85_result_delayed_u0=1'h0;
reg		reg_63b54bd2_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_6ca43d72_u0=1'h0;
reg		reg_2b115723_result_delayed_u0=1'h0;
reg		reg_45e011aa_result_delayed_u0=1'h0;
reg		reg_517738fd_result_delayed_result_delayed_u0=1'h0;
reg		reg_7a61a699_result_delayed_u0=1'h0;
reg		reg_4490a0a8_result_delayed_u0=1'h0;
reg		reg_25060cd9_u0=1'h0;
reg		reg_1dad4554_result_delayed_u0=1'h0;
reg		reg_6aa30297_result_delayed_u0=1'h0;
reg		reg_402ba1ce_u0=1'h0;
reg		reg_5325bac2_u0=1'h0;
reg		reg_53e492d4_result_delayed_u0=1'h0;
reg		reg_0d002d9e_result_delayed_u0=1'h0;
reg		reg_2927f9b8_result_delayed_u0=1'h0;
reg		reg_643841c9_u0=1'h0;
reg		reg_467e4f8d_u0=1'h0;
reg		reg_210fdd48_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_0c0741f4_u0=1'h0;
reg		reg_51727086_u0=1'h0;
reg		reg_015660ae_u0=1'h0;
reg		reg_6da5dd78_result_delayed_u0=1'h0;
reg		reg_07b4d1b4_u0=1'h0;
reg		reg_4ee47324_result_delayed_u0=1'h0;
reg		reg_457cf778_u0=1'h0;
reg		reg_5e114414_u0=1'h0;
reg		reg_68663660_u0=1'h0;
reg		reg_745b8e53_u0=1'h0;
reg		reg_75f2c8ed_result_delayed_u0=1'h0;
reg		reg_1aaa74b9_u0=1'h0;
reg		reg_4a513847_u0=1'h0;
reg		reg_068d86d5_result_delayed_result_delayed_u0=1'h0;
reg		reg_37e4d1fd_u0=1'h0;
reg		reg_123b2021_u0=1'h0;
reg		reg_37142796_result_delayed_u0=1'h0;
reg		reg_6b03bf9f_result_delayed_u0=1'h0;
reg		reg_2faca78c_result_delayed_result_delayed_u0=1'h0;
reg		reg_39988114_result_delayed_u0=1'h0;
reg		reg_0269f3e8_result_delayed_u0=1'h0;
reg		reg_3d184510_result_delayed_result_delayed_u0=1'h0;
reg		reg_4787c3ad_result_delayed_u0=1'h0;
reg		reg_393565d7_result_delayed_result_delayed_u0=1'h0;
reg		reg_330dd339_result_delayed_u0=1'h0;
reg		reg_61454769_u0=1'h0;
reg		reg_13d2c5ff_u0=1'h0;
reg		reg_3aa42c8a_u0=1'h0;
reg		reg_4a513847_result_delayed_u0=1'h0;
reg		reg_53436d73_u0=1'h0;
reg		reg_3d07ff30_u0=1'h0;
reg		reg_4302cd3b_u0=1'h0;
reg		reg_6fae0d94_u0=1'h0;
reg		reg_65238b18_u0=1'h0;
reg		reg_4d3f2823_result_delayed_u0=1'h0;
reg		reg_0269f3e8_result_delayed_result_delayed_u0=1'h0;
reg		reg_142e74f6_result_delayed_result_delayed_u0=1'h0;
reg		reg_1a329b29_result_delayed_u0=1'h0;
reg		reg_0dbaa983_result_delayed_result_delayed_u0=1'h0;
reg		reg_0848920e_u0=1'h0;
reg		reg_3027d020_result_delayed_u0=1'h0;
reg		reg_20dee699_u0=1'h0;
reg		reg_728c76f2_result_delayed_u0=1'h0;
reg		reg_5928537c_u0=1'h0;
reg		reg_6f4947f8_result_delayed_u0=1'h0;
reg		reg_6903fd17_result_delayed_result_delayed_u0=1'h0;
reg		reg_76680433_u0=1'h0;
reg		reg_643841c9_result_delayed_u0=1'h0;
reg		reg_170da16f_u0=1'h0;
reg		reg_63b54bd2_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_2b76cbc2_result_delayed_result_delayed_u0=1'h0;
reg		reg_07f782c9_result_delayed_u0=1'h0;
reg		reg_049c34f3_result_delayed_u0=1'h0;
reg		reg_19fcf5ae_result_delayed_u0=1'h0;
reg		reg_257da309_u0=1'h0;
reg		reg_550d08a9_result_delayed_u0=1'h0;
reg		reg_53915de4_u0=1'h0;
reg		reg_145a1005_result_delayed_u0=1'h0;
reg		reg_125f4827_u0=1'h0;
reg		reg_75f2c8ed_result_delayed_result_delayed_u0=1'h0;
reg		reg_20dee699_result_delayed_u0=1'h0;
reg		reg_660f9ef1_result_delayed_u0=1'h0;
reg		reg_3a3faffe_result_delayed_u0=1'h0;
reg		reg_37a25b06_result_delayed_u0=1'h0;
reg		reg_09925d27_result_delayed_u0=1'h0;
reg		reg_4beb2654_result_delayed_u0=1'h0;
wire		or_u1206_u0;
reg		reg_20fa067d_u0=1'h0;
reg		reg_57323713_result_delayed_result_delayed_u0=1'h0;
reg		reg_0d2097a9_u0=1'h0;
reg		reg_594f457a_result_delayed_result_delayed_u0=1'h0;
reg		reg_56f347a4_result_delayed_u0=1'h0;
reg		reg_2e9f4b96_result_delayed_u0=1'h0;
reg		reg_1aaa74b9_result_delayed_u0=1'h0;
reg		reg_0a6b2ffa_result_delayed_u0=1'h0;
reg		reg_20d7d0fd_result_delayed_u0=1'h0;
reg		reg_222a4f78_result_delayed_u0=1'h0;
reg		reg_0e961ae8_result_delayed_result_delayed_u0=1'h0;
reg		reg_417c43e2_u0=1'h0;
reg		reg_473d6b97_result_delayed_u0=1'h0;
reg		reg_11394f9b_u0=1'h0;
reg		reg_20703ad3_u0=1'h0;
reg		reg_0672d22b_result_delayed_u0=1'h0;
reg		reg_72fd2856_u0=1'h0;
reg		reg_0d2097a9_result_delayed_u0=1'h0;
reg		reg_23d37961_u0=1'h0;
reg		reg_7a53eec3_result_delayed_u0=1'h0;
reg		reg_41b4a953_result_delayed_u0=1'h0;
reg		reg_19be9d49_result_delayed_u0=1'h0;
reg		reg_1ae9a02b_u0=1'h0;
reg		reg_112873e3_u0=1'h0;
reg		reg_3cbd59f7_result_delayed_u0=1'h0;
reg		reg_4a513847_result_delayed_result_delayed_u0=1'h0;
reg		reg_745b8e53_result_delayed_u0=1'h0;
reg		reg_3e622eee_result_delayed_u0=1'h0;
reg		reg_47d47105_u0=1'h0;
reg		reg_47f58927_u0=1'h0;
reg		reg_73be9a15_result_delayed_u0=1'h0;
reg		reg_69dda494_result_delayed_u0=1'h0;
reg		reg_4fc71d19_u0=1'h0;
reg		reg_6cf4e62a_u0=1'h0;
reg		reg_20dee699_result_delayed_result_delayed_u0=1'h0;
reg		reg_79c318b3_result_delayed_u0=1'h0;
reg		reg_2eca9a1d_result_delayed_result_delayed_u0=1'h0;
reg		reg_2b115723_result_delayed_result_delayed_u0=1'h0;
reg		reg_45ddb9e8_result_delayed_u0=1'h0;
reg		reg_61454769_result_delayed_u0=1'h0;
reg		reg_7d2bf821_result_delayed_u0=1'h0;
reg		reg_112873e3_result_delayed_u0=1'h0;
reg		reg_7aa64abe_result_delayed_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_6ca43d72_result_delayed_u0=1'h0;
reg		reg_41b4a953_result_delayed_result_delayed_u0=1'h0;
reg		reg_3db89357_u0=1'h0;
reg		reg_1885f09c_result_delayed_result_delayed_u0=1'h0;
reg		reg_6535b053_result_delayed_u0=1'h0;
reg		reg_0a6b2ffa_result_delayed_result_delayed_u0=1'h0;
reg		reg_74b6d880_result_delayed_u0=1'h0;
reg		reg_4c652e93_u0=1'h0;
reg		reg_59d7b5da_result_delayed_u0=1'h0;
reg		reg_4b73b23b_result_delayed_u0=1'h0;
reg		reg_45f0eb0b_u0=1'h0;
reg		reg_7ad2c256_result_delayed_u0=1'h0;
reg		reg_2d74c675_u0=1'h0;
reg		reg_1aaa74b9_result_delayed_result_delayed_u0=1'h0;
reg		reg_67753870_u0=1'h0;
reg		reg_5ec29f05_result_delayed_u0=1'h0;
reg		reg_2376da04_result_delayed_u0=1'h0;
reg		reg_46627d70_u0=1'h0;
reg		reg_00ca0473_result_delayed_u0=1'h0;
reg		reg_741cf86b_result_delayed_result_delayed_u0=1'h0;
reg		reg_46861ff1_result_delayed_u0=1'h0;
reg		reg_45f0eb0b_result_delayed_u0=1'h0;
reg		reg_7ad2c256_result_delayed_result_delayed_u0=1'h0;
reg		reg_2e9f4b96_result_delayed_result_delayed_u0=1'h0;
reg		reg_0858480b_result_delayed_result_delayed_u0=1'h0;
reg		reg_4977a8c0_result_delayed_u0=1'h0;
reg		reg_1980ccbe_result_delayed_u0=1'h0;
reg		reg_3a57c6ba_result_delayed_u0=1'h0;
reg		reg_3b51abb4_result_delayed_u0=1'h0;
reg		reg_068d86d5_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_1a329b29_result_delayed_result_delayed_u0=1'h0;
reg		reg_2927f9b8_result_delayed_result_delayed_u0=1'h0;
reg		reg_794edd46_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_11bc6171_result_delayed_u0=1'h0;
reg		reg_45e011aa_result_delayed_result_delayed_u0=1'h0;
reg		reg_1f3d8a38_result_delayed_result_delayed_u0=1'h0;
reg		reg_45c4b9fe_result_delayed_result_delayed_u0=1'h0;
wire		and_u4068_u0;
reg		reg_19be9d49_result_delayed_result_delayed_u0=1'h0;
reg		reg_330dd339_result_delayed_result_delayed_u0=1'h0;
reg		reg_4f36662b_result_delayed_u0=1'h0;
reg		reg_41b4a953_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_29875567_result_delayed_result_delayed_u0=1'h0;
reg		reg_1b229062_u0=1'h0;
reg		reg_06c0f659_result_delayed_result_delayed_u0=1'h0;
reg		reg_10b12bf0_u0=1'h0;
reg		reg_7edc619f_u0=1'h0;
reg		reg_4ff7f3f0_result_delayed_u0=1'h0;
reg		reg_3027d020_result_delayed_result_delayed_u0=1'h0;
reg		reg_7e0c3547_u0=1'h0;
reg		reg_11bc6171_result_delayed_result_delayed_u0=1'h0;
reg		reg_41df9e8f_u0=1'h0;
reg		reg_3f89f30c_result_delayed_u0=1'h0;
reg		reg_46627d70_result_delayed_u0=1'h0;
reg		reg_7a53eec3_result_delayed_result_delayed_u0=1'h0;
reg		reg_3d07ff30_result_delayed_u0=1'h0;
reg		reg_45b236eb_u0=1'h0;
reg		reg_36d13294_result_delayed_u0=1'h0;
reg		reg_42c646a7_result_delayed_result_delayed_u0=1'h0;
reg		reg_45f0eb0b_result_delayed_result_delayed_u0=1'h0;
reg		and_delayed_u270=1'h0;
reg		reg_5e145a76_result_delayed_result_delayed_u0=1'h0;
reg		reg_2339dbf0_result_delayed_result_delayed_u0=1'h0;
reg		reg_4d562e3f_u0=1'h0;
reg		reg_3c50cd45_result_delayed_result_delayed_u0=1'h0;
reg		reg_6b2f3443_u0=1'h0;
reg		reg_6cf4e62a_result_delayed_u0=1'h0;
reg		reg_4274ae45_result_delayed_u0=1'h0;
reg		reg_4c652e93_result_delayed_u0=1'h0;
reg		reg_75f8153e_result_delayed_u0=1'h0;
reg		reg_53915de4_result_delayed_u0=1'h0;
reg		reg_1aaa74b9_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_07c27ed5_result_delayed_u0=1'h0;
reg		reg_4a513847_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_16604e6f_result_delayed_result_delayed_u0=1'h0;
reg		reg_6afd820d_result_delayed_u0=1'h0;
reg		reg_68663660_result_delayed_u0=1'h0;
reg		reg_0833f502_result_delayed_u0=1'h0;
reg		reg_4cae982d_result_delayed_result_delayed_u0=1'h0;
reg		reg_550541a9_result_delayed_u0=1'h0;
reg		reg_07b96631_result_delayed_u0=1'h0;
reg		reg_7e91f108_u0=1'h0;
reg		reg_358f4c1c_result_delayed_u0=1'h0;
reg		reg_6ceba0be_result_delayed_u0=1'h0;
reg		reg_7a61a699_result_delayed_result_delayed_u0=1'h0;
reg		reg_0848920e_result_delayed_u0=1'h0;
reg		reg_6b2f3443_result_delayed_u0=1'h0;
reg		reg_0d002d9e_result_delayed_result_delayed_u0=1'h0;
reg		reg_5325bac2_result_delayed_u0=1'h0;
reg		reg_2faca78c_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_4cbad8e5_result_delayed_result_delayed_u0=1'h0;
reg		reg_242dc5a0_result_delayed_u0=1'h0;
reg		reg_6abcb3ff_result_delayed_result_delayed_u0=1'h0;
reg		reg_48d7a190_result_delayed_u0=1'h0;
reg		reg_0e961ae8_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_1dad4554_result_delayed_result_delayed_u0=1'h0;
reg		reg_35c809c8_result_delayed_u0=1'h0;
reg		reg_1ae9a02b_result_delayed_u0=1'h0;
reg		reg_1aaa74b9_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_3726932e_result_delayed_u0=1'h0;
reg		reg_20d7d0fd_result_delayed_result_delayed_u0=1'h0;
reg		reg_29b64ddf_result_delayed_result_delayed_u0=1'h0;
reg		reg_125f4827_result_delayed_u0=1'h0;
reg		reg_79d4808b_result_delayed_result_delayed_u0=1'h0;
reg		reg_3c568577_result_delayed_u0=1'h0;
reg		reg_3aa42c8a_result_delayed_u0=1'h0;
reg		reg_16a5622b_result_delayed_u0=1'h0;
reg		reg_0120594a_result_delayed_u0=1'h0;
reg		reg_60829d18_result_delayed_u0=1'h0;
reg		reg_2eca9a1d_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_4c652e93_result_delayed_result_delayed_u0=1'h0;
reg		reg_21729149_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_4dc3c160_result_delayed_u0=1'h0;
reg		reg_2faca78c_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_14ea9829_result_delayed_u0=1'h0;
reg		reg_24743cb0_result_delayed_result_delayed_u0=1'h0;
reg		reg_20703ad3_result_delayed_u0=1'h0;
reg		reg_6b2f3443_result_delayed_result_delayed_u0=1'h0;
reg		reg_0e9d33d1_result_delayed_u0=1'h0;
reg		reg_330dd339_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_16a5622b_result_delayed_result_delayed_u0=1'h0;
reg		reg_63b54bd2_result_delayed_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_20d1a0f8_result_delayed_u0=1'h0;
reg		reg_2faca78c_result_delayed_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_20fa067d_result_delayed_u0=1'h0;
reg		reg_44c1644a_result_delayed_u0=1'h0;
reg		reg_23129694_result_delayed_u0=1'h0;
reg		reg_244f643a_result_delayed_u0=1'h0;
reg		reg_015660ae_result_delayed_u0=1'h0;
reg		reg_2eca9a1d_result_delayed_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_395b58c5_result_delayed_u0=1'h0;
reg		reg_5a3ed760_result_delayed_u0=1'h0;
reg		reg_0269f3e8_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_6b2f3443_result_delayed_result_delayed_result_delayed_u0=1'h0;
reg		reg_5f191bcf_u0=1'h0;
reg		reg_34efc738_u0=1'h0;
wire		and_u4069_u0;
wire		or_u1207_u0;
reg		reg_293a43e0_u0=1'h0;
wire		mux_u405_u0;
wire		or_u1208_u0;
reg		reg_3367383c_u0=1'h0;
wire		or_u1209_u0;
wire	[31:0]	mux_u406_u0;
reg		reg_5f191bcf_result_delayed_u0=1'h0;
wire		and_u4070_u0;
reg		reg_56c22f29_u0=1'h0;
reg		reg_3367383c_result_delayed_u0=1'h0;
reg		reg_56c22f29_result_delayed_u0=1'h0;
reg		reg_5f191bcf_result_delayed_result_delayed_u0=1'h0;
wire		or_u1210_u0;
wire		or_u1211_u0;
wire		or_u1212_u0;
wire		or_u1213_u0;
wire		and_u4071_u0;
wire		and_u4072_u0;
reg		and_delayed_u271_u0=1'h0;
wire signed	[31:0]	equals_u214_a_signed;
wire		equals_u214;
wire signed	[31:0]	equals_u214_b_signed;
wire		and_u4073_u0;
wire		and_u4074_u0;
wire		not_u649_u0;
wire		and_u4075_u0;
wire		not_u650_u0;
wire		and_u4076_u0;
wire signed	[31:0]	lessThan_u99_b_signed;
wire		lessThan_u99;
wire signed	[31:0]	lessThan_u99_a_signed;
wire		not_u651_u0;
wire		and_u4077_u0;
wire		and_u4078_u0;
wire		not_u652_u0;
wire		and_u4079_u0;
wire		and_u4080_u0;
wire	[31:0]	add;
wire		and_u4081_u0;
wire	[15:0]	simplePinWrite_u568;
wire		simplePinWrite_u569;
wire	[15:0]	simplePinWrite_u570;
wire	[31:0]	add_u575;
reg	[15:0]	syncEnable_u803=16'h0;
wire		and_u4082_u0;
wire	[15:0]	mux_u407_u0;
wire		and_u4083_u0;
reg		and_delayed_u272_u0=1'h0;
reg	[15:0]	syncEnable_u804_u0=16'h0;
reg		and_delayed_u273_u0=1'h0;
reg	[15:0]	syncEnable_u805_u0=16'h0;
wire	[15:0]	mux_u408_u0;
reg		reg_7f8418ac_u0=1'h0;
wire		and_u4084_u0;
reg	[31:0]	syncEnable_u806_u0=32'h0;
wire	[31:0]	mux_u409_u0;
wire		and_u4085_u0;
reg		and_delayed_u274_u0=1'h0;
wire		and_u4086_u0;
reg		and_delayed_u275_u0=1'h0;
reg	[15:0]	syncEnable_u807_u0=16'h0;
wire	[31:0]	mux_u410_u0;
reg		reg_79a785f7_u0=1'h0;
wire		and_u4087_u0;
wire	[15:0]	mux_u411_u0;
reg	[31:0]	syncEnable_u808_u0=32'h0;
wire		and_u4088_u0;
wire	[31:0]	mux_u412_u0;
wire		and_u4089_u0;
reg		and_delayed_u276_u0=1'h0;
reg	[31:0]	syncEnable_u809_u0=32'h0;
wire	[15:0]	mux_u413_u0;
reg		and_delayed_u277_u0=1'h0;
reg	[15:0]	syncEnable_u810_u0=16'h0;
wire		or_u1214_u0;
wire		mux_u414_u0;
reg	[31:0]	latch_7563f172_reg=32'h0;
wire	[31:0]	latch_7563f172_out;
wire	[15:0]	latch_4c497753_out;
reg	[15:0]	latch_4c497753_reg=16'h0;
wire		mux_u415_u0;
wire		or_u1215_u0;
reg		block_GO_delayed_u13=1'h0;
wire	[31:0]	mux_u416_u0;
wire		or_u1216_u0;
wire		or_u1217_u0;
wire	[31:0]	mux_u417_u0;
wire		and_u4090_u0;
wire	[15:0]	mux_u418_u0;
wire		or_u1218_u0;
wire	[31:0]	mux_u419_u0;
reg	[15:0]	fbReg_Out1Portvalue_u5=16'h0;
reg	[31:0]	fbReg_temp_fsmOldState_resized_LH3_xy_8_u0=32'h0;
reg		syncEnable_u811_u0=1'h0;
reg		loopControl_u10=1'h0;
wire	[31:0]	mux_u420_u0;
wire		or_u1219_u0;
wire		or_u1220_u0;
reg		reg_4dbfab2c_u0=1'h0;
wire		or_u1221_u0;
wire	[31:0]	mux_u421_u0;
wire		mux_u422_u0;
wire		or_u1222_u0;
wire		or_u1223_u0;
wire		mux_u423_u0;
reg		reg_585ee52a_u0=1'h0;
assign lessThan_a_unsigned=port_1bba0a1c_;
assign lessThan_b_unsigned=16'h40;
assign lessThan=lessThan_a_unsigned<lessThan_b_unsigned;
assign equals_a_unsigned=port_1bba0a1c_;
assign equals_b_unsigned=16'h40;
assign equals=equals_a_unsigned==equals_b_unsigned;
assign lessThan_u98_a_unsigned=port_4c65738f_;
assign lessThan_u98_b_unsigned=16'h8;
assign lessThan_u98=lessThan_u98_a_unsigned<lessThan_u98_b_unsigned;
assign andOp=equals&lessThan_u98;
assign equals_u212_a_unsigned=port_4c65738f_;
assign equals_u212_b_unsigned=16'h8;
assign equals_u212=equals_u212_a_unsigned==equals_u212_b_unsigned;
assign equals_u213_a_signed={31'b0, port_6cb7d4b7_};
assign equals_u213_b_signed=32'h0;
assign equals_u213=equals_u213_a_signed==equals_u213_b_signed;
assign not_u645_u0=~equals_u213;
assign and_u4058_u0=and_u4090_u0&equals_u213;
assign and_u4059_u0=and_u4090_u0&not_u645_u0;
assign andOp_u213=lessThan&port_157e6b5b_;
assign and_u4060_u0=and_u4071_u0&not_u646_u0;
assign not_u646_u0=~andOp_u213;
assign and_u4061_u0=and_u4071_u0&andOp_u213;
assign simplePinWrite=and_u4070_u0&{1{and_u4070_u0}};
assign not_u647_u0=~andOp;
assign and_u4062_u0=and_u4069_u0&andOp;
assign and_u4063_u0=and_u4069_u0&not_u647_u0;
assign simplePinWrite_u566=and_u4067_u0&{1{and_u4067_u0}};
assign and_u4064_u0=and_u4068_u0&not_u648_u0;
assign not_u648_u0=~equals_u212;
assign and_u4065_u0=and_u4068_u0&equals_u212;
assign simplePinWrite_u567=and_u4066_u0&{1{and_u4066_u0}};
assign and_u4066_u0=and_u4065_u0&and_u4068_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4985bd85_u0<=1'h0;
else reg_4985bd85_u0<=reg_6b924716_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_35c809c8_u0<=1'h0;
else reg_35c809c8_u0<=reg_67e7177f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5760cf63_u0<=1'h0;
else reg_5760cf63_u0<=reg_343be065_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6fb08fb4_u0<=1'h0;
else reg_6fb08fb4_u0<=reg_3c7ba446_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4ff7f3f0_u0<=1'h0;
else reg_4ff7f3f0_u0<=reg_2cb66d26_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3027d020_u0<=1'h0;
else reg_3027d020_u0<=reg_0c0741f4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_794edd46_u0<=1'h0;
else reg_794edd46_u0<=reg_745b8e53_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3726932e_u0<=1'h0;
else reg_3726932e_u0<=reg_1a329b29_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3d184510_u0<=1'h0;
else reg_3d184510_u0<=reg_3c0ef12e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_59d7b5da_u0<=1'h0;
else reg_59d7b5da_u0<=reg_45c4b9fe_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_16604e6f_u0<=1'h0;
else reg_16604e6f_u0<=reg_512aac58_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6903fd17_u0<=1'h0;
else reg_6903fd17_u0<=reg_11394f9b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7aa64abe_u0<=1'h0;
else reg_7aa64abe_u0<=reg_2b115723_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1885f09c_u0<=1'h0;
else reg_1885f09c_u0<=reg_4ee47324_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2faca78c_u0<=1'h0;
else reg_2faca78c_u0<=reg_794edd46_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_57323713_u0<=1'h0;
else reg_57323713_u0<=reg_19be9d49_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_20d1a0f8_u0<=1'h0;
else reg_20d1a0f8_u0<=reg_413e1dbb_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_20d7d0fd_u0<=1'h0;
else reg_20d7d0fd_u0<=reg_746c5835_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4787c3ad_u0<=1'h0;
else reg_4787c3ad_u0<=reg_49a5b9d0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4274ae45_u0<=1'h0;
else reg_4274ae45_u0<=reg_69c13d7a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2b115723_u0<=1'h0;
else reg_2b115723_u0<=reg_2d8038cc_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_330dd339_u0<=1'h0;
else reg_330dd339_u0<=reg_16a5622b_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6aa30297_u0<=1'h0;
else reg_6aa30297_u0<=reg_3c50cd45_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_45ddb9e8_u0<=1'h0;
else reg_45ddb9e8_u0<=reg_257da309_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_594f457a_u0<=1'h0;
else reg_594f457a_u0<=reg_4b73b23b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_74b6d880_u0<=1'h0;
else reg_74b6d880_u0<=reg_21f11516_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4490a0a8_u0<=1'h0;
else reg_4490a0a8_u0<=reg_7bcb7712_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3cb65c8f_u0<=1'h0;
else reg_3cb65c8f_u0<=reg_2d178d82_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0dbaa983_u0<=1'h0;
else reg_0dbaa983_u0<=reg_4beb2654_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_45c4b9fe_u0<=1'h0;
else reg_45c4b9fe_u0<=reg_671babf3_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_21729149_u0<=1'h0;
else reg_21729149_u0<=reg_6d8fa179_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3c7ba446_u0<=1'h0;
else reg_3c7ba446_u0<=reg_3cb65c8f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1b5e971f_u0<=1'h0;
else reg_1b5e971f_u0<=reg_0c1a90ca_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_36d13294_u0<=1'h0;
else reg_36d13294_u0<=reg_3d3b0167_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_210fdd48_u0<=1'h0;
else reg_210fdd48_u0<=reg_393565d7_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_45e011aa_u0<=1'h0;
else reg_45e011aa_u0<=reg_3cbd59f7_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_21729149_result_delayed_u0<=1'h0;
else reg_21729149_result_delayed_u0<=reg_21729149_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_55e64da9_u0<=1'h0;
else reg_55e64da9_u0<=reg_309c310d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_19fcf5ae_u0<=1'h0;
else reg_19fcf5ae_u0<=reg_618a90a2_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0858480b_u0<=1'h0;
else reg_0858480b_u0<=reg_4f36662b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_21729149_result_delayed_result_delayed_u0<=1'h0;
else reg_21729149_result_delayed_result_delayed_u0<=reg_21729149_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6ceba0be_u0<=1'h0;
else reg_6ceba0be_u0<=reg_7edc619f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_068d86d5_u0<=1'h0;
else reg_068d86d5_u0<=reg_550d08a9_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_746c5835_u0<=1'h0;
else reg_746c5835_u0<=reg_238aead6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0672d22b_u0<=1'h0;
else reg_0672d22b_u0<=reg_55e64da9_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3d3b0167_u0<=1'h0;
else reg_3d3b0167_u0<=reg_6af44a24_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_55e64da9_result_delayed_u0<=1'h0;
else reg_55e64da9_result_delayed_u0<=reg_55e64da9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_343be065_u0<=1'h0;
else reg_343be065_u0<=reg_39988114_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_145a1005_u0<=1'h0;
else reg_145a1005_u0<=reg_1b229062_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4cbad8e5_u0<=1'h0;
else reg_4cbad8e5_u0<=reg_145a1005_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_42c646a7_u0<=1'h0;
else reg_42c646a7_u0<=reg_2a0b1f83_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5e145a76_u0<=1'h0;
else reg_5e145a76_u0<=reg_53436d73_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_63b54bd2_u0<=1'h0;
else reg_63b54bd2_u0<=reg_123b2021_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_29b64ddf_u0<=1'h0;
else reg_29b64ddf_u0<=reg_36d13294_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0120594a_u0<=1'h0;
else reg_0120594a_u0<=reg_741cf86b_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_049c34f3_u0<=1'h0;
else reg_049c34f3_u0<=reg_50958802_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_244f643a_u0<=1'h0;
else reg_244f643a_u0<=reg_5f70cbfe_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_49a5b9d0_u0<=1'h0;
else reg_49a5b9d0_u0<=reg_594f457a_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_741cf86b_u0<=1'h0;
else reg_741cf86b_u0<=reg_29875567_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0e961ae8_u0<=1'h0;
else reg_0e961ae8_u0<=reg_0833f502_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_728c76f2_u0<=1'h0;
else reg_728c76f2_u0<=reg_660f9ef1_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0e961ae8_result_delayed_u0<=1'h0;
else reg_0e961ae8_result_delayed_u0<=reg_0e961ae8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_37142796_u0<=1'h0;
else reg_37142796_u0<=reg_45e011aa_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4cae982d_u0<=1'h0;
else reg_4cae982d_u0<=reg_457cf778_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6b924716_u0<=1'h0;
else reg_6b924716_u0<=reg_14042498_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7ad2c256_u0<=1'h0;
else reg_7ad2c256_u0<=reg_37142796_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_413e1dbb_u0<=1'h0;
else reg_413e1dbb_u0<=reg_4787c3ad_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3f89f30c_u0<=1'h0;
else reg_3f89f30c_u0<=reg_51727086_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_44c1644a_u0<=1'h0;
else reg_44c1644a_u0<=reg_6aa9532f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3e622eee_u0<=1'h0;
else reg_3e622eee_u0<=reg_7a61a699_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_39988114_u0<=1'h0;
else reg_39988114_u0<=reg_2339dbf0_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_16a5622b_u0<=1'h0;
else reg_16a5622b_u0<=reg_4c652e93_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5f70cbfe_u0<=1'h0;
else reg_5f70cbfe_u0<=reg_3a57c6ba_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a53eec3_u0<=1'h0;
else reg_7a53eec3_u0<=reg_1dad4554_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2d178d82_u0<=1'h0;
else reg_2d178d82_u0<=reg_2f1102bc_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_50958802_u0<=1'h0;
else reg_50958802_u0<=reg_01dd2487_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_430f0398_u0<=1'h0;
else reg_430f0398_u0<=reg_5091b5e2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_67e7177f_u0<=1'h0;
else reg_67e7177f_u0<=reg_4a3d5eec_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_06c0f659_u0<=1'h0;
else reg_06c0f659_u0<=reg_20dee699_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_210fdd48_result_delayed_u0<=1'h0;
else reg_210fdd48_result_delayed_u0<=reg_210fdd48_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_14042498_u0<=1'h0;
else reg_14042498_u0<=reg_75f8153e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6b03bf9f_u0<=1'h0;
else reg_6b03bf9f_u0<=reg_3c568577_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7e53b6cf_u0<=1'h0;
else reg_7e53b6cf_u0<=and_u4068_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0d002d9e_u0<=1'h0;
else reg_0d002d9e_u0<=reg_07f782c9_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2927f9b8_u0<=1'h0;
else reg_2927f9b8_u0<=reg_222a4f78_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4dc3c160_u0<=1'h0;
else reg_4dc3c160_u0<=reg_64d83df2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_37a25b06_u0<=1'h0;
else reg_37a25b06_u0<=reg_7213e342_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_473d6b97_u0<=1'h0;
else reg_473d6b97_u0<=reg_72fd2856_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_068d86d5_result_delayed_u0<=1'h0;
else reg_068d86d5_result_delayed_u0<=reg_068d86d5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_550541a9_u0<=1'h0;
else reg_550541a9_u0<=reg_22e61fae_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3131c19c_u0<=1'h0;
else reg_3131c19c_u0<=reg_06c0f659_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6f4947f8_u0<=1'h0;
else reg_6f4947f8_u0<=reg_53e492d4_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_16604e6f_result_delayed_u0<=1'h0;
else reg_16604e6f_result_delayed_u0<=reg_16604e6f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2b76cbc2_u0<=1'h0;
else reg_2b76cbc2_u0<=reg_45b236eb_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_09925d27_u0<=1'h0;
else reg_09925d27_u0<=reg_430f0398_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00ca0473_u0<=1'h0;
else reg_00ca0473_u0<=reg_5928537c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_63b54bd2_result_delayed_u0<=1'h0;
else reg_63b54bd2_result_delayed_u0<=reg_63b54bd2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_69c13d7a_u0<=1'h0;
else reg_69c13d7a_u0<=reg_74b6d880_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5f70cbfe_result_delayed_u0<=1'h0;
else reg_5f70cbfe_result_delayed_u0<=reg_5f70cbfe_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_14ea9829_u0<=1'h0;
else reg_14ea9829_u0<=reg_41df9e8f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_24743cb0_u0<=1'h0;
else reg_24743cb0_u0<=reg_07c27ed5_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_75f8153e_u0<=1'h0;
else reg_75f8153e_u0<=reg_4a513847_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6b924716_result_delayed_u0<=1'h0;
else reg_6b924716_result_delayed_u0<=reg_6b924716_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2339dbf0_u0<=1'h0;
else reg_2339dbf0_u0<=reg_2927f9b8_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_11bc6171_u0<=1'h0;
else reg_11bc6171_u0<=reg_1f3d8a38_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6af44a24_u0<=1'h0;
else reg_6af44a24_u0<=reg_37f5df2f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0c1a90ca_u0<=1'h0;
else reg_0c1a90ca_u0<=reg_330dd339_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4a3d5eec_u0<=1'h0;
else reg_4a3d5eec_u0<=reg_142e74f6_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2339dbf0_result_delayed_u0<=1'h0;
else reg_2339dbf0_result_delayed_u0<=reg_2339dbf0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_29b64ddf_result_delayed_u0<=1'h0;
else reg_29b64ddf_result_delayed_u0<=reg_29b64ddf_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0858480b_result_delayed_u0<=1'h0;
else reg_0858480b_result_delayed_u0<=reg_0858480b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2eca9a1d_u0<=1'h0;
else reg_2eca9a1d_u0<=reg_5e114414_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_142e74f6_u0<=1'h0;
else reg_142e74f6_u0<=reg_3fe03efe_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7bcb7712_u0<=1'h0;
else reg_7bcb7712_u0<=reg_4fc71d19_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_37f5df2f_u0<=1'h0;
else reg_37f5df2f_u0<=reg_6d25a062_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2b76cbc2_result_delayed_u0<=1'h0;
else reg_2b76cbc2_result_delayed_u0<=reg_2b76cbc2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6da5dd78_u0<=1'h0;
else reg_6da5dd78_u0<=reg_35c809c8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_794edd46_result_delayed_u0<=1'h0;
else reg_794edd46_result_delayed_u0<=reg_794edd46_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_29875567_u0<=1'h0;
else reg_29875567_u0<=reg_24743cb0_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_55e64da9_result_delayed_result_delayed_u0<=1'h0;
else reg_55e64da9_result_delayed_result_delayed_u0<=reg_55e64da9_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_393565d7_u0<=1'h0;
else reg_393565d7_u0<=reg_395b58c5_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3b51abb4_u0<=1'h0;
else reg_3b51abb4_u0<=reg_76680433_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_21f11516_u0<=1'h0;
else reg_21f11516_u0<=reg_3a5d4aa0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_41b4a953_u0<=1'h0;
else reg_41b4a953_u0<=reg_53915de4_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_671babf3_u0<=1'h0;
else reg_671babf3_u0<=reg_44c1644a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3a57c6ba_u0<=1'h0;
else reg_3a57c6ba_u0<=reg_6f4947f8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6afd820d_u0<=1'h0;
else reg_6afd820d_u0<=reg_45f0eb0b_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_393565d7_result_delayed_u0<=1'h0;
else reg_393565d7_result_delayed_u0<=reg_393565d7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6d8fa179_u0<=1'h0;
else reg_6d8fa179_u0<=reg_3d184510_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_19be9d49_u0<=1'h0;
else reg_19be9d49_u0<=reg_4cbad8e5_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a61a699_u0<=1'h0;
else reg_7a61a699_u0<=reg_07b4d1b4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1dad4554_u0<=1'h0;
else reg_1dad4554_u0<=reg_473d6b97_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3a5d4aa0_u0<=1'h0;
else reg_3a5d4aa0_u0<=reg_467e4f8d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_660f9ef1_u0<=1'h0;
else reg_660f9ef1_u0<=reg_57323713_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1f3d8a38_u0<=1'h0;
else reg_1f3d8a38_u0<=reg_42c646a7_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_430f0398_result_delayed_u0<=1'h0;
else reg_430f0398_result_delayed_u0<=reg_430f0398_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7aa64abe_result_delayed_u0<=1'h0;
else reg_7aa64abe_result_delayed_u0<=reg_7aa64abe_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_210fdd48_result_delayed_result_delayed_u0<=1'h0;
else reg_210fdd48_result_delayed_result_delayed_u0<=reg_210fdd48_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2e9f4b96_u0<=1'h0;
else reg_2e9f4b96_u0<=reg_7a53eec3_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7d2bf821_u0<=1'h0;
else reg_7d2bf821_u0<=reg_5760cf63_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5760cf63_result_delayed_u0<=1'h0;
else reg_5760cf63_result_delayed_u0<=reg_5760cf63_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2eca9a1d_result_delayed_u0<=1'h0;
else reg_2eca9a1d_result_delayed_u0<=reg_2eca9a1d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3c50cd45_u0<=1'h0;
else reg_3c50cd45_u0<=reg_6b03bf9f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4cae982d_result_delayed_u0<=1'h0;
else reg_4cae982d_result_delayed_u0<=reg_4cae982d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_07c27ed5_u0<=1'h0;
else reg_07c27ed5_u0<=reg_21729149_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1f3d8a38_result_delayed_u0<=1'h0;
else reg_1f3d8a38_result_delayed_u0<=reg_1f3d8a38_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1a329b29_u0<=1'h0;
else reg_1a329b29_u0<=reg_5a3ed760_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4d3f2823_u0<=1'h0;
else reg_4d3f2823_u0<=reg_7ad08748_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4f36662b_u0<=1'h0;
else reg_4f36662b_u0<=reg_6535b053_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3fe03efe_u0<=1'h0;
else reg_3fe03efe_u0<=reg_20703ad3_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_75f2c8ed_u0<=1'h0;
else reg_75f2c8ed_u0<=reg_28ebf99a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3c0ef12e_u0<=1'h0;
else reg_3c0ef12e_u0<=reg_068d86d5_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3c568577_u0<=1'h0;
else reg_3c568577_u0<=reg_529137a1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1885f09c_result_delayed_u0<=1'h0;
else reg_1885f09c_result_delayed_u0<=reg_1885f09c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2c201504_u0<=1'h0;
else reg_2c201504_u0<=reg_37a25b06_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_618a90a2_u0<=1'h0;
else reg_618a90a2_u0<=reg_3726932e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5e145a76_result_delayed_u0<=1'h0;
else reg_5e145a76_result_delayed_u0<=reg_5e145a76_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_618a90a2_result_delayed_u0<=1'h0;
else reg_618a90a2_result_delayed_u0<=reg_618a90a2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_64d83df2_u0<=1'h0;
else reg_64d83df2_u0<=reg_4d3f2823_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_594f457a_result_delayed_u0<=1'h0;
else reg_594f457a_result_delayed_u0<=reg_594f457a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7aa64abe_result_delayed_result_delayed_u0<=1'h0;
else reg_7aa64abe_result_delayed_result_delayed_u0<=reg_7aa64abe_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_529137a1_u0<=1'h0;
else reg_529137a1_u0<=reg_79c318b3_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_53e492d4_u0<=1'h0;
else reg_53e492d4_u0<=reg_2c201504_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0833f502_u0<=1'h0;
else reg_0833f502_u0<=reg_3131c19c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1b5e971f_result_delayed_u0<=1'h0;
else reg_1b5e971f_result_delayed_u0<=reg_1b5e971f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0c1a90ca_result_delayed_u0<=1'h0;
else reg_0c1a90ca_result_delayed_u0<=reg_0c1a90ca_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_142e74f6_result_delayed_u0<=1'h0;
else reg_142e74f6_result_delayed_u0<=reg_142e74f6_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_07f782c9_u0<=1'h0;
else reg_07f782c9_u0<=reg_049c34f3_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1980ccbe_u0<=1'h0;
else reg_1980ccbe_u0<=reg_6da5dd78_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_63b54bd2_result_delayed_result_delayed_u0<=1'h0;
else reg_63b54bd2_result_delayed_result_delayed_u0<=reg_63b54bd2_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_45c4b9fe_result_delayed_u0<=1'h0;
else reg_45c4b9fe_result_delayed_u0<=reg_45c4b9fe_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3d3b0167_result_delayed_u0<=1'h0;
else reg_3d3b0167_result_delayed_u0<=reg_3d3b0167_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6af44a24_result_delayed_u0<=1'h0;
else reg_6af44a24_result_delayed_u0<=reg_6af44a24_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6abcb3ff_u0<=1'h0;
else reg_6abcb3ff_u0<=reg_75f2c8ed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6d25a062_u0<=1'h0;
else reg_6d25a062_u0<=reg_23129694_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_48d7a190_u0<=1'h0;
else reg_48d7a190_u0<=reg_37e4d1fd_u0;
end
assign mux_u404=(and_u4067_u0)?1'h1:1'h0;
assign or_u1205_u0=and_u4067_u0|and_u4066_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4b73b23b_u0<=1'h0;
else reg_4b73b23b_u0<=reg_003f51b2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_22e61fae_u0<=1'h0;
else reg_22e61fae_u0<=reg_3f89f30c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_69dda494_u0<=1'h0;
else reg_69dda494_u0<=reg_320deb94_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3cbd59f7_u0<=1'h0;
else reg_3cbd59f7_u0<=reg_6ca43d72_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0e9d33d1_u0<=1'h0;
else reg_0e9d33d1_u0<=reg_14ea9829_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2d8038cc_u0<=1'h0;
else reg_2d8038cc_u0<=reg_13d2c5ff_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7213e342_u0<=1'h0;
else reg_7213e342_u0<=reg_7aa64abe_result_delayed_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_222a4f78_u0<=1'h0;
else reg_222a4f78_u0<=reg_4dc3c160_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0dbaa983_result_delayed_u0<=1'h0;
else reg_0dbaa983_result_delayed_u0<=reg_0dbaa983_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3c50cd45_result_delayed_u0<=1'h0;
else reg_3c50cd45_result_delayed_u0<=reg_3c50cd45_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_56f347a4_u0<=1'h0;
else reg_56f347a4_u0<=reg_20d1a0f8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01dd2487_u0<=1'h0;
else reg_01dd2487_u0<=and_delayed_u270;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_238aead6_u0<=1'h0;
else reg_238aead6_u0<=reg_6fb08fb4_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5a3ed760_u0<=1'h0;
else reg_5a3ed760_u0<=reg_47f58927_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_79d4808b_u0<=1'h0;
else reg_79d4808b_u0<=reg_1aaa74b9_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6fb08fb4_result_delayed_u0<=1'h0;
else reg_6fb08fb4_result_delayed_u0<=reg_6fb08fb4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3d184510_result_delayed_u0<=1'h0;
else reg_3d184510_result_delayed_u0<=reg_3d184510_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_430f0398_result_delayed_result_delayed_u0<=1'h0;
else reg_430f0398_result_delayed_result_delayed_u0<=reg_430f0398_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6535b053_u0<=1'h0;
else reg_6535b053_u0<=reg_3b51abb4_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7aa64abe_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_7aa64abe_result_delayed_result_delayed_result_delayed_u0<=reg_7aa64abe_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6d25a062_result_delayed_u0<=1'h0;
else reg_6d25a062_result_delayed_u0<=reg_6d25a062_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_618a90a2_result_delayed_result_delayed_u0<=1'h0;
else reg_618a90a2_result_delayed_result_delayed_u0<=reg_618a90a2_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_79c318b3_u0<=1'h0;
else reg_79c318b3_u0<=reg_4985bd85_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_28ebf99a_u0<=1'h0;
else reg_28ebf99a_u0<=reg_1b5e971f_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2376da04_u0<=1'h0;
else reg_2376da04_u0<=reg_6aa30297_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_512aac58_u0<=1'h0;
else reg_512aac58_u0<=reg_25060cd9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5091b5e2_u0<=1'h0;
else reg_5091b5e2_u0<=reg_56f347a4_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_741cf86b_result_delayed_u0<=1'h0;
else reg_741cf86b_result_delayed_u0<=reg_741cf86b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6abcb3ff_result_delayed_u0<=1'h0;
else reg_6abcb3ff_result_delayed_u0<=reg_6abcb3ff_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_46861ff1_u0<=1'h0;
else reg_46861ff1_u0<=reg_0dbaa983_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3131c19c_result_delayed_u0<=1'h0;
else reg_3131c19c_result_delayed_u0<=reg_3131c19c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0269f3e8_u0<=1'h0;
else reg_0269f3e8_u0<=reg_5325bac2_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1b5e971f_result_delayed_result_delayed_u0<=1'h0;
else reg_1b5e971f_result_delayed_result_delayed_u0<=reg_1b5e971f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_23129694_u0<=1'h0;
else reg_23129694_u0<=reg_7101c0a1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6aa9532f_u0<=1'h0;
else reg_6aa9532f_u0<=reg_19fcf5ae_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2a0b1f83_u0<=1'h0;
else reg_2a0b1f83_u0<=reg_222c2bb3_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_07b96631_u0<=1'h0;
else reg_07b96631_u0<=reg_65238b18_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_517738fd_u0<=1'h0;
else reg_517738fd_u0<=reg_4490a0a8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_42c646a7_result_delayed_u0<=1'h0;
else reg_42c646a7_result_delayed_u0<=reg_42c646a7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01dd2487_result_delayed_u0<=1'h0;
else reg_01dd2487_result_delayed_u0<=reg_01dd2487_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_242dc5a0_u0<=1'h0;
else reg_242dc5a0_u0<=reg_16604e6f_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_003f51b2_u0<=1'h0;
else reg_003f51b2_u0<=reg_2b76cbc2_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2cb66d26_u0<=1'h0;
else reg_2cb66d26_u0<=reg_517738fd_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_794edd46_result_delayed_result_delayed_u0<=1'h0;
else reg_794edd46_result_delayed_result_delayed_u0<=reg_794edd46_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_309c310d_u0<=1'h0;
else reg_309c310d_u0<=reg_5ec29f05_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0a6b2ffa_u0<=1'h0;
else reg_0a6b2ffa_u0<=reg_0d2097a9_result_delayed_u0;
end
assign and_u4067_u0=and_u4062_u0&and_u4069_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_517738fd_result_delayed_u0<=1'h0;
else reg_517738fd_result_delayed_u0<=reg_517738fd_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_358f4c1c_u0<=1'h0;
else reg_358f4c1c_u0<=reg_7d2bf821_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7ad08748_u0<=1'h0;
else reg_7ad08748_u0<=reg_3027d020_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_320deb94_u0<=1'h0;
else reg_320deb94_u0<=reg_59d7b5da_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_60829d18_u0<=1'h0;
else reg_60829d18_u0<=reg_0858480b_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_395b58c5_u0<=1'h0;
else reg_395b58c5_u0<=reg_170da16f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_222c2bb3_u0<=1'h0;
else reg_222c2bb3_u0<=reg_67753870_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_57323713_result_delayed_u0<=1'h0;
else reg_57323713_result_delayed_u0<=reg_57323713_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7101c0a1_u0<=1'h0;
else reg_7101c0a1_u0<=reg_0d002d9e_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_550d08a9_u0<=1'h0;
else reg_550d08a9_u0<=reg_2e9f4b96_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6903fd17_result_delayed_u0<=1'h0;
else reg_6903fd17_result_delayed_u0<=reg_6903fd17_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2faca78c_result_delayed_u0<=1'h0;
else reg_2faca78c_result_delayed_u0<=reg_2faca78c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_343be065_result_delayed_u0<=1'h0;
else reg_343be065_result_delayed_u0<=reg_343be065_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_73be9a15_u0<=1'h0;
else reg_73be9a15_u0<=reg_29b64ddf_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7213e342_result_delayed_u0<=1'h0;
else reg_7213e342_result_delayed_u0<=reg_7213e342_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2f1102bc_u0<=1'h0;
else reg_2f1102bc_u0<=reg_2d74c675_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3cb65c8f_result_delayed_u0<=1'h0;
else reg_3cb65c8f_result_delayed_u0<=reg_3cb65c8f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7aa64abe_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_7aa64abe_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_7aa64abe_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4977a8c0_u0<=1'h0;
else reg_4977a8c0_u0<=reg_0e9d33d1_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2c201504_result_delayed_u0<=1'h0;
else reg_2c201504_result_delayed_u0<=reg_2c201504_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4cbad8e5_result_delayed_u0<=1'h0;
else reg_4cbad8e5_result_delayed_u0<=reg_4cbad8e5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_06c0f659_result_delayed_u0<=1'h0;
else reg_06c0f659_result_delayed_u0<=reg_06c0f659_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6d8fa179_result_delayed_u0<=1'h0;
else reg_6d8fa179_result_delayed_u0<=reg_6d8fa179_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_29875567_result_delayed_u0<=1'h0;
else reg_29875567_result_delayed_u0<=reg_29875567_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4beb2654_u0<=1'h0;
else reg_4beb2654_u0<=reg_0a6b2ffa_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4ee47324_u0<=1'h0;
else reg_4ee47324_u0<=reg_210fdd48_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3a3faffe_u0<=1'h0;
else reg_3a3faffe_u0<=reg_402ba1ce_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_79d4808b_result_delayed_u0<=1'h0;
else reg_79d4808b_result_delayed_u0<=reg_79d4808b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_24743cb0_result_delayed_u0<=1'h0;
else reg_24743cb0_result_delayed_u0<=reg_24743cb0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_343be065_result_delayed_result_delayed_u0<=1'h0;
else reg_343be065_result_delayed_result_delayed_u0<=reg_343be065_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5ec29f05_u0<=1'h0;
else reg_5ec29f05_u0<=reg_07b96631_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4985bd85_result_delayed_u0<=1'h0;
else reg_4985bd85_result_delayed_u0<=reg_4985bd85_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_63b54bd2_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_63b54bd2_result_delayed_result_delayed_result_delayed_u0<=reg_63b54bd2_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6ca43d72_u0<=1'h0;
else reg_6ca43d72_u0<=reg_45ddb9e8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2b115723_result_delayed_u0<=1'h0;
else reg_2b115723_result_delayed_u0<=reg_2b115723_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_45e011aa_result_delayed_u0<=1'h0;
else reg_45e011aa_result_delayed_u0<=reg_45e011aa_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_517738fd_result_delayed_result_delayed_u0<=1'h0;
else reg_517738fd_result_delayed_result_delayed_u0<=reg_517738fd_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a61a699_result_delayed_u0<=1'h0;
else reg_7a61a699_result_delayed_u0<=reg_7a61a699_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4490a0a8_result_delayed_u0<=1'h0;
else reg_4490a0a8_result_delayed_u0<=reg_4490a0a8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_25060cd9_u0<=1'h0;
else reg_25060cd9_u0<=reg_69dda494_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1dad4554_result_delayed_u0<=1'h0;
else reg_1dad4554_result_delayed_u0<=reg_1dad4554_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6aa30297_result_delayed_u0<=1'h0;
else reg_6aa30297_result_delayed_u0<=reg_6aa30297_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_402ba1ce_u0<=1'h0;
else reg_402ba1ce_u0<=reg_09925d27_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5325bac2_u0<=1'h0;
else reg_5325bac2_u0<=reg_4d562e3f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_53e492d4_result_delayed_u0<=1'h0;
else reg_53e492d4_result_delayed_u0<=reg_53e492d4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0d002d9e_result_delayed_u0<=1'h0;
else reg_0d002d9e_result_delayed_u0<=reg_0d002d9e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2927f9b8_result_delayed_u0<=1'h0;
else reg_2927f9b8_result_delayed_u0<=reg_2927f9b8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_643841c9_u0<=1'h0;
else reg_643841c9_u0<=reg_6abcb3ff_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_467e4f8d_u0<=1'h0;
else reg_467e4f8d_u0<=reg_2376da04_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_210fdd48_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_210fdd48_result_delayed_result_delayed_result_delayed_u0<=reg_210fdd48_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0c0741f4_u0<=1'h0;
else reg_0c0741f4_u0<=reg_1885f09c_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_51727086_u0<=1'h0;
else reg_51727086_u0<=reg_728c76f2_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_015660ae_u0<=1'h0;
else reg_015660ae_u0<=reg_4302cd3b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6da5dd78_result_delayed_u0<=1'h0;
else reg_6da5dd78_result_delayed_u0<=reg_6da5dd78_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_07b4d1b4_u0<=1'h0;
else reg_07b4d1b4_u0<=reg_3db89357_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4ee47324_result_delayed_u0<=1'h0;
else reg_4ee47324_result_delayed_u0<=reg_4ee47324_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_457cf778_u0<=1'h0;
else reg_457cf778_u0<=reg_41b4a953_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5e114414_u0<=1'h0;
else reg_5e114414_u0<=reg_242dc5a0_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_68663660_u0<=1'h0;
else reg_68663660_u0<=reg_2eca9a1d_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_745b8e53_u0<=1'h0;
else reg_745b8e53_u0<=reg_6b2f3443_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_75f2c8ed_result_delayed_u0<=1'h0;
else reg_75f2c8ed_result_delayed_u0<=reg_75f2c8ed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1aaa74b9_u0<=1'h0;
else reg_1aaa74b9_u0<=reg_643841c9_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4a513847_u0<=1'h0;
else reg_4a513847_u0<=reg_6fae0d94_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_068d86d5_result_delayed_result_delayed_u0<=1'h0;
else reg_068d86d5_result_delayed_result_delayed_u0<=reg_068d86d5_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_37e4d1fd_u0<=1'h0;
else reg_37e4d1fd_u0<=reg_0269f3e8_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_123b2021_u0<=1'h0;
else reg_123b2021_u0<=reg_6903fd17_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_37142796_result_delayed_u0<=1'h0;
else reg_37142796_result_delayed_u0<=reg_37142796_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6b03bf9f_result_delayed_u0<=1'h0;
else reg_6b03bf9f_result_delayed_u0<=reg_6b03bf9f_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2faca78c_result_delayed_result_delayed_u0<=1'h0;
else reg_2faca78c_result_delayed_result_delayed_u0<=reg_2faca78c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_39988114_result_delayed_u0<=1'h0;
else reg_39988114_result_delayed_u0<=reg_39988114_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0269f3e8_result_delayed_u0<=1'h0;
else reg_0269f3e8_result_delayed_u0<=reg_0269f3e8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3d184510_result_delayed_result_delayed_u0<=1'h0;
else reg_3d184510_result_delayed_result_delayed_u0<=reg_3d184510_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4787c3ad_result_delayed_u0<=1'h0;
else reg_4787c3ad_result_delayed_u0<=reg_4787c3ad_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_393565d7_result_delayed_result_delayed_u0<=1'h0;
else reg_393565d7_result_delayed_result_delayed_u0<=reg_393565d7_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_330dd339_result_delayed_u0<=1'h0;
else reg_330dd339_result_delayed_u0<=reg_330dd339_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_61454769_u0<=1'h0;
else reg_61454769_u0<=reg_46861ff1_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_13d2c5ff_u0<=1'h0;
else reg_13d2c5ff_u0<=reg_68663660_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3aa42c8a_u0<=1'h0;
else reg_3aa42c8a_u0<=reg_48d7a190_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4a513847_result_delayed_u0<=1'h0;
else reg_4a513847_result_delayed_u0<=reg_4a513847_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_53436d73_u0<=1'h0;
else reg_53436d73_u0<=reg_3a3faffe_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3d07ff30_u0<=1'h0;
else reg_3d07ff30_u0<=reg_3e622eee_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4302cd3b_u0<=1'h0;
else reg_4302cd3b_u0<=reg_244f643a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6fae0d94_u0<=1'h0;
else reg_6fae0d94_u0<=reg_417c43e2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_65238b18_u0<=1'h0;
else reg_65238b18_u0<=reg_7ad2c256_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4d3f2823_result_delayed_u0<=1'h0;
else reg_4d3f2823_result_delayed_u0<=reg_4d3f2823_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0269f3e8_result_delayed_result_delayed_u0<=1'h0;
else reg_0269f3e8_result_delayed_result_delayed_u0<=reg_0269f3e8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_142e74f6_result_delayed_result_delayed_u0<=1'h0;
else reg_142e74f6_result_delayed_result_delayed_u0<=reg_142e74f6_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1a329b29_result_delayed_u0<=1'h0;
else reg_1a329b29_result_delayed_u0<=reg_1a329b29_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0dbaa983_result_delayed_result_delayed_u0<=1'h0;
else reg_0dbaa983_result_delayed_result_delayed_u0<=reg_0dbaa983_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0848920e_u0<=1'h0;
else reg_0848920e_u0<=reg_015660ae_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3027d020_result_delayed_u0<=1'h0;
else reg_3027d020_result_delayed_u0<=reg_3027d020_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_20dee699_u0<=1'h0;
else reg_20dee699_u0<=reg_63b54bd2_result_delayed_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_728c76f2_result_delayed_u0<=1'h0;
else reg_728c76f2_result_delayed_u0<=reg_728c76f2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5928537c_u0<=1'h0;
else reg_5928537c_u0<=reg_23d37961_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6f4947f8_result_delayed_u0<=1'h0;
else reg_6f4947f8_result_delayed_u0<=reg_6f4947f8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6903fd17_result_delayed_result_delayed_u0<=1'h0;
else reg_6903fd17_result_delayed_result_delayed_u0<=reg_6903fd17_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_76680433_u0<=1'h0;
else reg_76680433_u0<=reg_5e145a76_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_643841c9_result_delayed_u0<=1'h0;
else reg_643841c9_result_delayed_u0<=reg_643841c9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_170da16f_u0<=1'h0;
else reg_170da16f_u0<=reg_0672d22b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_63b54bd2_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_63b54bd2_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_63b54bd2_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2b76cbc2_result_delayed_result_delayed_u0<=1'h0;
else reg_2b76cbc2_result_delayed_result_delayed_u0<=reg_2b76cbc2_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_07f782c9_result_delayed_u0<=1'h0;
else reg_07f782c9_result_delayed_u0<=reg_07f782c9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_049c34f3_result_delayed_u0<=1'h0;
else reg_049c34f3_result_delayed_u0<=reg_049c34f3_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_19fcf5ae_result_delayed_u0<=1'h0;
else reg_19fcf5ae_result_delayed_u0<=reg_19fcf5ae_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_257da309_u0<=1'h0;
else reg_257da309_u0<=reg_0120594a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_550d08a9_result_delayed_u0<=1'h0;
else reg_550d08a9_result_delayed_u0<=reg_550d08a9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_53915de4_u0<=1'h0;
else reg_53915de4_u0<=reg_61454769_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_145a1005_result_delayed_u0<=1'h0;
else reg_145a1005_result_delayed_u0<=reg_145a1005_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_125f4827_u0<=1'h0;
else reg_125f4827_u0<=reg_4ff7f3f0_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_75f2c8ed_result_delayed_result_delayed_u0<=1'h0;
else reg_75f2c8ed_result_delayed_result_delayed_u0<=reg_75f2c8ed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_20dee699_result_delayed_u0<=1'h0;
else reg_20dee699_result_delayed_u0<=reg_20dee699_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_660f9ef1_result_delayed_u0<=1'h0;
else reg_660f9ef1_result_delayed_u0<=reg_660f9ef1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3a3faffe_result_delayed_u0<=1'h0;
else reg_3a3faffe_result_delayed_u0<=reg_3a3faffe_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_37a25b06_result_delayed_u0<=1'h0;
else reg_37a25b06_result_delayed_u0<=reg_37a25b06_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_09925d27_result_delayed_u0<=1'h0;
else reg_09925d27_result_delayed_u0<=reg_09925d27_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4beb2654_result_delayed_u0<=1'h0;
else reg_4beb2654_result_delayed_u0<=reg_4beb2654_u0;
end
assign or_u1206_u0=reg_550541a9_result_delayed_u0|reg_7e53b6cf_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_20fa067d_u0<=1'h0;
else reg_20fa067d_u0<=reg_7e91f108_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_57323713_result_delayed_result_delayed_u0<=1'h0;
else reg_57323713_result_delayed_result_delayed_u0<=reg_57323713_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0d2097a9_u0<=1'h0;
else reg_0d2097a9_u0<=reg_20fa067d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_594f457a_result_delayed_result_delayed_u0<=1'h0;
else reg_594f457a_result_delayed_result_delayed_u0<=reg_594f457a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_56f347a4_result_delayed_u0<=1'h0;
else reg_56f347a4_result_delayed_u0<=reg_56f347a4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2e9f4b96_result_delayed_u0<=1'h0;
else reg_2e9f4b96_result_delayed_u0<=reg_2e9f4b96_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1aaa74b9_result_delayed_u0<=1'h0;
else reg_1aaa74b9_result_delayed_u0<=reg_1aaa74b9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0a6b2ffa_result_delayed_u0<=1'h0;
else reg_0a6b2ffa_result_delayed_u0<=reg_0a6b2ffa_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_20d7d0fd_result_delayed_u0<=1'h0;
else reg_20d7d0fd_result_delayed_u0<=reg_20d7d0fd_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_222a4f78_result_delayed_u0<=1'h0;
else reg_222a4f78_result_delayed_u0<=reg_222a4f78_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0e961ae8_result_delayed_result_delayed_u0<=1'h0;
else reg_0e961ae8_result_delayed_result_delayed_u0<=reg_0e961ae8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_417c43e2_u0<=1'h0;
else reg_417c43e2_u0<=reg_4977a8c0_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_473d6b97_result_delayed_u0<=1'h0;
else reg_473d6b97_result_delayed_u0<=reg_473d6b97_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_11394f9b_u0<=1'h0;
else reg_11394f9b_u0<=reg_73be9a15_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_20703ad3_u0<=1'h0;
else reg_20703ad3_u0<=reg_3d07ff30_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0672d22b_result_delayed_u0<=1'h0;
else reg_0672d22b_result_delayed_u0<=reg_0672d22b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_72fd2856_u0<=1'h0;
else reg_72fd2856_u0<=reg_0848920e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0d2097a9_result_delayed_u0<=1'h0;
else reg_0d2097a9_result_delayed_u0<=reg_0d2097a9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_23d37961_u0<=1'h0;
else reg_23d37961_u0<=reg_1980ccbe_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a53eec3_result_delayed_u0<=1'h0;
else reg_7a53eec3_result_delayed_u0<=reg_7a53eec3_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_41b4a953_result_delayed_u0<=1'h0;
else reg_41b4a953_result_delayed_u0<=reg_41b4a953_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_19be9d49_result_delayed_u0<=1'h0;
else reg_19be9d49_result_delayed_u0<=reg_19be9d49_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1ae9a02b_u0<=1'h0;
else reg_1ae9a02b_u0<=reg_3aa42c8a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_112873e3_u0<=1'h0;
else reg_112873e3_u0<=reg_47d47105_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3cbd59f7_result_delayed_u0<=1'h0;
else reg_3cbd59f7_result_delayed_u0<=reg_3cbd59f7_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4a513847_result_delayed_result_delayed_u0<=1'h0;
else reg_4a513847_result_delayed_result_delayed_u0<=reg_4a513847_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_745b8e53_result_delayed_u0<=1'h0;
else reg_745b8e53_result_delayed_u0<=reg_745b8e53_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3e622eee_result_delayed_u0<=1'h0;
else reg_3e622eee_result_delayed_u0<=reg_3e622eee_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_47d47105_u0<=1'h0;
else reg_47d47105_u0<=reg_46627d70_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_47f58927_u0<=1'h0;
else reg_47f58927_u0<=reg_112873e3_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_73be9a15_result_delayed_u0<=1'h0;
else reg_73be9a15_result_delayed_u0<=reg_73be9a15_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_69dda494_result_delayed_u0<=1'h0;
else reg_69dda494_result_delayed_u0<=reg_69dda494_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4fc71d19_u0<=1'h0;
else reg_4fc71d19_u0<=reg_11bc6171_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6cf4e62a_u0<=1'h0;
else reg_6cf4e62a_u0<=reg_10b12bf0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_20dee699_result_delayed_result_delayed_u0<=1'h0;
else reg_20dee699_result_delayed_result_delayed_u0<=reg_20dee699_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_79c318b3_result_delayed_u0<=1'h0;
else reg_79c318b3_result_delayed_u0<=reg_79c318b3_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2eca9a1d_result_delayed_result_delayed_u0<=1'h0;
else reg_2eca9a1d_result_delayed_result_delayed_u0<=reg_2eca9a1d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2b115723_result_delayed_result_delayed_u0<=1'h0;
else reg_2b115723_result_delayed_result_delayed_u0<=reg_2b115723_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_45ddb9e8_result_delayed_u0<=1'h0;
else reg_45ddb9e8_result_delayed_u0<=reg_45ddb9e8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_61454769_result_delayed_u0<=1'h0;
else reg_61454769_result_delayed_u0<=reg_61454769_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7d2bf821_result_delayed_u0<=1'h0;
else reg_7d2bf821_result_delayed_u0<=reg_7d2bf821_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_112873e3_result_delayed_u0<=1'h0;
else reg_112873e3_result_delayed_u0<=reg_112873e3_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7aa64abe_result_delayed_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_7aa64abe_result_delayed_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_7aa64abe_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6ca43d72_result_delayed_u0<=1'h0;
else reg_6ca43d72_result_delayed_u0<=reg_6ca43d72_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_41b4a953_result_delayed_result_delayed_u0<=1'h0;
else reg_41b4a953_result_delayed_result_delayed_u0<=reg_41b4a953_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3db89357_u0<=1'h0;
else reg_3db89357_u0<=reg_7e0c3547_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1885f09c_result_delayed_result_delayed_u0<=1'h0;
else reg_1885f09c_result_delayed_result_delayed_u0<=reg_1885f09c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6535b053_result_delayed_u0<=1'h0;
else reg_6535b053_result_delayed_u0<=reg_6535b053_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0a6b2ffa_result_delayed_result_delayed_u0<=1'h0;
else reg_0a6b2ffa_result_delayed_result_delayed_u0<=reg_0a6b2ffa_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_74b6d880_result_delayed_u0<=1'h0;
else reg_74b6d880_result_delayed_u0<=reg_74b6d880_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4c652e93_u0<=1'h0;
else reg_4c652e93_u0<=reg_6ceba0be_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_59d7b5da_result_delayed_u0<=1'h0;
else reg_59d7b5da_result_delayed_u0<=reg_59d7b5da_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4b73b23b_result_delayed_u0<=1'h0;
else reg_4b73b23b_result_delayed_u0<=reg_4b73b23b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_45f0eb0b_u0<=1'h0;
else reg_45f0eb0b_u0<=reg_2faca78c_result_delayed_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7ad2c256_result_delayed_u0<=1'h0;
else reg_7ad2c256_result_delayed_u0<=reg_7ad2c256_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2d74c675_u0<=1'h0;
else reg_2d74c675_u0<=reg_00ca0473_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1aaa74b9_result_delayed_result_delayed_u0<=1'h0;
else reg_1aaa74b9_result_delayed_result_delayed_u0<=reg_1aaa74b9_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_67753870_u0<=1'h0;
else reg_67753870_u0<=reg_4274ae45_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5ec29f05_result_delayed_u0<=1'h0;
else reg_5ec29f05_result_delayed_u0<=reg_5ec29f05_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2376da04_result_delayed_u0<=1'h0;
else reg_2376da04_result_delayed_u0<=reg_2376da04_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_46627d70_u0<=1'h0;
else reg_46627d70_u0<=reg_6afd820d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00ca0473_result_delayed_u0<=1'h0;
else reg_00ca0473_result_delayed_u0<=reg_00ca0473_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_741cf86b_result_delayed_result_delayed_u0<=1'h0;
else reg_741cf86b_result_delayed_result_delayed_u0<=reg_741cf86b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_46861ff1_result_delayed_u0<=1'h0;
else reg_46861ff1_result_delayed_u0<=reg_46861ff1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_45f0eb0b_result_delayed_u0<=1'h0;
else reg_45f0eb0b_result_delayed_u0<=reg_45f0eb0b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7ad2c256_result_delayed_result_delayed_u0<=1'h0;
else reg_7ad2c256_result_delayed_result_delayed_u0<=reg_7ad2c256_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2e9f4b96_result_delayed_result_delayed_u0<=1'h0;
else reg_2e9f4b96_result_delayed_result_delayed_u0<=reg_2e9f4b96_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0858480b_result_delayed_result_delayed_u0<=1'h0;
else reg_0858480b_result_delayed_result_delayed_u0<=reg_0858480b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4977a8c0_result_delayed_u0<=1'h0;
else reg_4977a8c0_result_delayed_u0<=reg_4977a8c0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1980ccbe_result_delayed_u0<=1'h0;
else reg_1980ccbe_result_delayed_u0<=reg_1980ccbe_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3a57c6ba_result_delayed_u0<=1'h0;
else reg_3a57c6ba_result_delayed_u0<=reg_3a57c6ba_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3b51abb4_result_delayed_u0<=1'h0;
else reg_3b51abb4_result_delayed_u0<=reg_3b51abb4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_068d86d5_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_068d86d5_result_delayed_result_delayed_result_delayed_u0<=reg_068d86d5_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1a329b29_result_delayed_result_delayed_u0<=1'h0;
else reg_1a329b29_result_delayed_result_delayed_u0<=reg_1a329b29_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2927f9b8_result_delayed_result_delayed_u0<=1'h0;
else reg_2927f9b8_result_delayed_result_delayed_u0<=reg_2927f9b8_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_794edd46_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_794edd46_result_delayed_result_delayed_result_delayed_u0<=reg_794edd46_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_11bc6171_result_delayed_u0<=1'h0;
else reg_11bc6171_result_delayed_u0<=reg_11bc6171_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_45e011aa_result_delayed_result_delayed_u0<=1'h0;
else reg_45e011aa_result_delayed_result_delayed_u0<=reg_45e011aa_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1f3d8a38_result_delayed_result_delayed_u0<=1'h0;
else reg_1f3d8a38_result_delayed_result_delayed_u0<=reg_1f3d8a38_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_45c4b9fe_result_delayed_result_delayed_u0<=1'h0;
else reg_45c4b9fe_result_delayed_result_delayed_u0<=reg_45c4b9fe_result_delayed_u0;
end
assign and_u4068_u0=and_u4063_u0&and_u4069_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_19be9d49_result_delayed_result_delayed_u0<=1'h0;
else reg_19be9d49_result_delayed_result_delayed_u0<=reg_19be9d49_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_330dd339_result_delayed_result_delayed_u0<=1'h0;
else reg_330dd339_result_delayed_result_delayed_u0<=reg_330dd339_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4f36662b_result_delayed_u0<=1'h0;
else reg_4f36662b_result_delayed_u0<=reg_4f36662b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_41b4a953_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_41b4a953_result_delayed_result_delayed_result_delayed_u0<=reg_41b4a953_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_29875567_result_delayed_result_delayed_u0<=1'h0;
else reg_29875567_result_delayed_result_delayed_u0<=reg_29875567_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1b229062_u0<=1'h0;
else reg_1b229062_u0<=reg_4cae982d_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_06c0f659_result_delayed_result_delayed_u0<=1'h0;
else reg_06c0f659_result_delayed_result_delayed_u0<=reg_06c0f659_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_10b12bf0_u0<=1'h0;
else reg_10b12bf0_u0<=reg_125f4827_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7edc619f_u0<=1'h0;
else reg_7edc619f_u0<=reg_0e961ae8_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4ff7f3f0_result_delayed_u0<=1'h0;
else reg_4ff7f3f0_result_delayed_u0<=reg_4ff7f3f0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3027d020_result_delayed_result_delayed_u0<=1'h0;
else reg_3027d020_result_delayed_result_delayed_u0<=reg_3027d020_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7e0c3547_u0<=1'h0;
else reg_7e0c3547_u0<=reg_6cf4e62a_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_11bc6171_result_delayed_result_delayed_u0<=1'h0;
else reg_11bc6171_result_delayed_result_delayed_u0<=reg_11bc6171_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_41df9e8f_u0<=1'h0;
else reg_41df9e8f_u0<=reg_79d4808b_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3f89f30c_result_delayed_u0<=1'h0;
else reg_3f89f30c_result_delayed_u0<=reg_3f89f30c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_46627d70_result_delayed_u0<=1'h0;
else reg_46627d70_result_delayed_u0<=reg_46627d70_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a53eec3_result_delayed_result_delayed_u0<=1'h0;
else reg_7a53eec3_result_delayed_result_delayed_u0<=reg_7a53eec3_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3d07ff30_result_delayed_u0<=1'h0;
else reg_3d07ff30_result_delayed_u0<=reg_3d07ff30_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_45b236eb_u0<=1'h0;
else reg_45b236eb_u0<=reg_358f4c1c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_36d13294_result_delayed_u0<=1'h0;
else reg_36d13294_result_delayed_u0<=reg_36d13294_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_42c646a7_result_delayed_result_delayed_u0<=1'h0;
else reg_42c646a7_result_delayed_result_delayed_u0<=reg_42c646a7_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_45f0eb0b_result_delayed_result_delayed_u0<=1'h0;
else reg_45f0eb0b_result_delayed_result_delayed_u0<=reg_45f0eb0b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u270<=1'h0;
else and_delayed_u270<=and_u4067_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5e145a76_result_delayed_result_delayed_u0<=1'h0;
else reg_5e145a76_result_delayed_result_delayed_u0<=reg_5e145a76_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2339dbf0_result_delayed_result_delayed_u0<=1'h0;
else reg_2339dbf0_result_delayed_result_delayed_u0<=reg_2339dbf0_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4d562e3f_u0<=1'h0;
else reg_4d562e3f_u0<=reg_60829d18_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3c50cd45_result_delayed_result_delayed_u0<=1'h0;
else reg_3c50cd45_result_delayed_result_delayed_u0<=reg_3c50cd45_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6b2f3443_u0<=1'h0;
else reg_6b2f3443_u0<=reg_20d7d0fd_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6cf4e62a_result_delayed_u0<=1'h0;
else reg_6cf4e62a_result_delayed_u0<=reg_6cf4e62a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4274ae45_result_delayed_u0<=1'h0;
else reg_4274ae45_result_delayed_u0<=reg_4274ae45_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4c652e93_result_delayed_u0<=1'h0;
else reg_4c652e93_result_delayed_u0<=reg_4c652e93_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_75f8153e_result_delayed_u0<=1'h0;
else reg_75f8153e_result_delayed_u0<=reg_75f8153e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_53915de4_result_delayed_u0<=1'h0;
else reg_53915de4_result_delayed_u0<=reg_53915de4_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1aaa74b9_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_1aaa74b9_result_delayed_result_delayed_result_delayed_u0<=reg_1aaa74b9_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_07c27ed5_result_delayed_u0<=1'h0;
else reg_07c27ed5_result_delayed_u0<=reg_07c27ed5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4a513847_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_4a513847_result_delayed_result_delayed_result_delayed_u0<=reg_4a513847_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_16604e6f_result_delayed_result_delayed_u0<=1'h0;
else reg_16604e6f_result_delayed_result_delayed_u0<=reg_16604e6f_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6afd820d_result_delayed_u0<=1'h0;
else reg_6afd820d_result_delayed_u0<=reg_6afd820d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_68663660_result_delayed_u0<=1'h0;
else reg_68663660_result_delayed_u0<=reg_68663660_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0833f502_result_delayed_u0<=1'h0;
else reg_0833f502_result_delayed_u0<=reg_0833f502_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4cae982d_result_delayed_result_delayed_u0<=1'h0;
else reg_4cae982d_result_delayed_result_delayed_u0<=reg_4cae982d_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_550541a9_result_delayed_u0<=1'h0;
else reg_550541a9_result_delayed_u0<=reg_550541a9_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_07b96631_result_delayed_u0<=1'h0;
else reg_07b96631_result_delayed_u0<=reg_07b96631_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7e91f108_u0<=1'h0;
else reg_7e91f108_u0<=reg_1ae9a02b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_358f4c1c_result_delayed_u0<=1'h0;
else reg_358f4c1c_result_delayed_u0<=reg_358f4c1c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6ceba0be_result_delayed_u0<=1'h0;
else reg_6ceba0be_result_delayed_u0<=reg_6ceba0be_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7a61a699_result_delayed_result_delayed_u0<=1'h0;
else reg_7a61a699_result_delayed_result_delayed_u0<=reg_7a61a699_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0848920e_result_delayed_u0<=1'h0;
else reg_0848920e_result_delayed_u0<=reg_0848920e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6b2f3443_result_delayed_u0<=1'h0;
else reg_6b2f3443_result_delayed_u0<=reg_6b2f3443_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0d002d9e_result_delayed_result_delayed_u0<=1'h0;
else reg_0d002d9e_result_delayed_result_delayed_u0<=reg_0d002d9e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5325bac2_result_delayed_u0<=1'h0;
else reg_5325bac2_result_delayed_u0<=reg_5325bac2_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2faca78c_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_2faca78c_result_delayed_result_delayed_result_delayed_u0<=reg_2faca78c_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4cbad8e5_result_delayed_result_delayed_u0<=1'h0;
else reg_4cbad8e5_result_delayed_result_delayed_u0<=reg_4cbad8e5_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_242dc5a0_result_delayed_u0<=1'h0;
else reg_242dc5a0_result_delayed_u0<=reg_242dc5a0_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6abcb3ff_result_delayed_result_delayed_u0<=1'h0;
else reg_6abcb3ff_result_delayed_result_delayed_u0<=reg_6abcb3ff_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_48d7a190_result_delayed_u0<=1'h0;
else reg_48d7a190_result_delayed_u0<=reg_48d7a190_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0e961ae8_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_0e961ae8_result_delayed_result_delayed_result_delayed_u0<=reg_0e961ae8_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1dad4554_result_delayed_result_delayed_u0<=1'h0;
else reg_1dad4554_result_delayed_result_delayed_u0<=reg_1dad4554_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_35c809c8_result_delayed_u0<=1'h0;
else reg_35c809c8_result_delayed_u0<=reg_35c809c8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1ae9a02b_result_delayed_u0<=1'h0;
else reg_1ae9a02b_result_delayed_u0<=reg_1ae9a02b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1aaa74b9_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_1aaa74b9_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_1aaa74b9_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3726932e_result_delayed_u0<=1'h0;
else reg_3726932e_result_delayed_u0<=reg_3726932e_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_20d7d0fd_result_delayed_result_delayed_u0<=1'h0;
else reg_20d7d0fd_result_delayed_result_delayed_u0<=reg_20d7d0fd_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_29b64ddf_result_delayed_result_delayed_u0<=1'h0;
else reg_29b64ddf_result_delayed_result_delayed_u0<=reg_29b64ddf_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_125f4827_result_delayed_u0<=1'h0;
else reg_125f4827_result_delayed_u0<=reg_125f4827_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_79d4808b_result_delayed_result_delayed_u0<=1'h0;
else reg_79d4808b_result_delayed_result_delayed_u0<=reg_79d4808b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3c568577_result_delayed_u0<=1'h0;
else reg_3c568577_result_delayed_u0<=reg_3c568577_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3aa42c8a_result_delayed_u0<=1'h0;
else reg_3aa42c8a_result_delayed_u0<=reg_3aa42c8a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_16a5622b_result_delayed_u0<=1'h0;
else reg_16a5622b_result_delayed_u0<=reg_16a5622b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0120594a_result_delayed_u0<=1'h0;
else reg_0120594a_result_delayed_u0<=reg_0120594a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_60829d18_result_delayed_u0<=1'h0;
else reg_60829d18_result_delayed_u0<=reg_60829d18_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2eca9a1d_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_2eca9a1d_result_delayed_result_delayed_result_delayed_u0<=reg_2eca9a1d_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4c652e93_result_delayed_result_delayed_u0<=1'h0;
else reg_4c652e93_result_delayed_result_delayed_u0<=reg_4c652e93_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_21729149_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_21729149_result_delayed_result_delayed_result_delayed_u0<=reg_21729149_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4dc3c160_result_delayed_u0<=1'h0;
else reg_4dc3c160_result_delayed_u0<=reg_4dc3c160_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2faca78c_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_2faca78c_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_2faca78c_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_14ea9829_result_delayed_u0<=1'h0;
else reg_14ea9829_result_delayed_u0<=reg_14ea9829_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_24743cb0_result_delayed_result_delayed_u0<=1'h0;
else reg_24743cb0_result_delayed_result_delayed_u0<=reg_24743cb0_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_20703ad3_result_delayed_u0<=1'h0;
else reg_20703ad3_result_delayed_u0<=reg_20703ad3_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6b2f3443_result_delayed_result_delayed_u0<=1'h0;
else reg_6b2f3443_result_delayed_result_delayed_u0<=reg_6b2f3443_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0e9d33d1_result_delayed_u0<=1'h0;
else reg_0e9d33d1_result_delayed_u0<=reg_0e9d33d1_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_330dd339_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_330dd339_result_delayed_result_delayed_result_delayed_u0<=reg_330dd339_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_16a5622b_result_delayed_result_delayed_u0<=1'h0;
else reg_16a5622b_result_delayed_result_delayed_u0<=reg_16a5622b_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_63b54bd2_result_delayed_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_63b54bd2_result_delayed_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_63b54bd2_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_20d1a0f8_result_delayed_u0<=1'h0;
else reg_20d1a0f8_result_delayed_u0<=reg_20d1a0f8_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2faca78c_result_delayed_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_2faca78c_result_delayed_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_2faca78c_result_delayed_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_20fa067d_result_delayed_u0<=1'h0;
else reg_20fa067d_result_delayed_u0<=reg_20fa067d_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_44c1644a_result_delayed_u0<=1'h0;
else reg_44c1644a_result_delayed_u0<=reg_44c1644a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_23129694_result_delayed_u0<=1'h0;
else reg_23129694_result_delayed_u0<=reg_23129694_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_244f643a_result_delayed_u0<=1'h0;
else reg_244f643a_result_delayed_u0<=reg_244f643a_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_015660ae_result_delayed_u0<=1'h0;
else reg_015660ae_result_delayed_u0<=reg_015660ae_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_2eca9a1d_result_delayed_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_2eca9a1d_result_delayed_result_delayed_result_delayed_result_delayed_u0<=reg_2eca9a1d_result_delayed_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_395b58c5_result_delayed_u0<=1'h0;
else reg_395b58c5_result_delayed_u0<=reg_395b58c5_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5a3ed760_result_delayed_u0<=1'h0;
else reg_5a3ed760_result_delayed_u0<=reg_5a3ed760_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0269f3e8_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_0269f3e8_result_delayed_result_delayed_result_delayed_u0<=reg_0269f3e8_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6b2f3443_result_delayed_result_delayed_result_delayed_u0<=1'h0;
else reg_6b2f3443_result_delayed_result_delayed_result_delayed_u0<=reg_6b2f3443_result_delayed_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5f191bcf_u0<=1'h0;
else reg_5f191bcf_u0<=and_u4070_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_34efc738_u0<=1'h0;
else reg_34efc738_u0<=reg_293a43e0_u0;
end
assign and_u4069_u0=and_u4060_u0&and_u4071_u0;
assign or_u1207_u0=and_u4070_u0|and_u4067_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_293a43e0_u0<=1'h0;
else reg_293a43e0_u0<=reg_56c22f29_result_delayed_u0;
end
assign mux_u405_u0=(and_u4070_u0)?1'h1:mux_u404;
assign or_u1208_u0=and_u4070_u0|or_u1205_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3367383c_u0<=1'h0;
else reg_3367383c_u0<=reg_5f191bcf_result_delayed_result_delayed_u0;
end
assign or_u1209_u0=and_u4070_u0|and_u4067_u0;
assign mux_u406_u0=(and_u4070_u0)?32'h8:32'h200;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5f191bcf_result_delayed_u0<=1'h0;
else reg_5f191bcf_result_delayed_u0<=reg_5f191bcf_u0;
end
assign and_u4070_u0=and_u4061_u0&and_u4071_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_56c22f29_u0<=1'h0;
else reg_56c22f29_u0<=reg_3367383c_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_3367383c_result_delayed_u0<=1'h0;
else reg_3367383c_result_delayed_u0<=reg_3367383c_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_56c22f29_result_delayed_u0<=1'h0;
else reg_56c22f29_result_delayed_u0<=reg_56c22f29_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_5f191bcf_result_delayed_result_delayed_u0<=1'h0;
else reg_5f191bcf_result_delayed_result_delayed_u0<=reg_5f191bcf_result_delayed_u0;
end
assign or_u1210_u0=and_u4070_u0|and_u4067_u0;
assign or_u1211_u0=reg_34efc738_u0|or_u1206_u0;
assign or_u1212_u0=and_u4070_u0|and_u4067_u0;
assign or_u1213_u0=or_u1211_u0|and_delayed_u271_u0;
assign and_u4071_u0=and_u4058_u0&and_u4090_u0;
assign and_u4072_u0=and_u4059_u0&and_u4090_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u271_u0<=1'h0;
else and_delayed_u271_u0<=and_u4072_u0;
end
assign equals_u214_a_signed={31'b0, port_6cb7d4b7_};
assign equals_u214_b_signed=32'h1;
assign equals_u214=equals_u214_a_signed==equals_u214_b_signed;
assign and_u4073_u0=and_u4090_u0&equals_u214;
assign and_u4074_u0=and_u4090_u0&not_u649_u0;
assign not_u649_u0=~equals_u214;
assign and_u4075_u0=and_u4089_u0&port_202620a3_;
assign not_u650_u0=~port_202620a3_;
assign and_u4076_u0=and_u4089_u0&not_u650_u0;
assign lessThan_u99_a_signed=port_639e94f2_;
assign lessThan_u99_b_signed=port_072ed7ee_;
assign lessThan_u99=lessThan_u99_a_signed<lessThan_u99_b_signed;
assign not_u651_u0=~lessThan_u99;
assign and_u4077_u0=and_u4087_u0&not_u651_u0;
assign and_u4078_u0=and_u4087_u0&lessThan_u99;
assign not_u652_u0=~port_7fb2b3af_;
assign and_u4079_u0=and_u4085_u0&port_7fb2b3af_;
assign and_u4080_u0=and_u4085_u0&not_u652_u0;
assign add=port_639e94f2_+32'h0;
assign and_u4081_u0=and_u4082_u0&port_03915889_;
assign simplePinWrite_u568=16'h1&{16{1'h1}};
assign simplePinWrite_u569=and_u4082_u0&{1{and_u4082_u0}};
assign simplePinWrite_u570=port_5c53ee9c_;
assign add_u575=port_639e94f2_+32'h1;
always @(posedge CLK)
begin
if (and_u4082_u0)
syncEnable_u803<=port_5c53ee9c_;
end
assign and_u4082_u0=and_u4079_u0&and_u4085_u0;
assign mux_u407_u0=(and_delayed_u272_u0)?syncEnable_u803:syncEnable_u804_u0;
assign and_u4083_u0=and_u4080_u0&and_u4085_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u272_u0<=1'h0;
else and_delayed_u272_u0<=and_u4082_u0;
end
always @(posedge CLK)
begin
if (and_u4085_u0)
syncEnable_u804_u0<=mux_u418_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u273_u0<=1'h0;
else and_delayed_u273_u0<=and_u4083_u0;
end
always @(posedge CLK)
begin
if (and_u4087_u0)
syncEnable_u805_u0<=mux_u418_u0;
end
assign mux_u408_u0=(reg_7f8418ac_u0)?syncEnable_u805_u0:mux_u407_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_7f8418ac_u0<=1'h0;
else reg_7f8418ac_u0<=and_u4084_u0;
end
assign and_u4084_u0=and_u4077_u0&and_u4087_u0;
always @(posedge CLK)
begin
if (and_u4087_u0)
syncEnable_u806_u0<=mux_u419_u0;
end
assign mux_u409_u0=(reg_7f8418ac_u0)?32'h0:syncEnable_u806_u0;
assign and_u4085_u0=and_u4078_u0&and_u4087_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u274_u0<=1'h0;
else and_delayed_u274_u0<=and_u4085_u0;
end
assign and_u4086_u0=and_u4076_u0&and_u4089_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u275_u0<=1'h0;
else and_delayed_u275_u0<=and_u4086_u0;
end
always @(posedge CLK)
begin
if (and_u4089_u0)
syncEnable_u807_u0<=mux_u418_u0;
end
assign mux_u410_u0=(reg_79a785f7_u0)?mux_u409_u0:syncEnable_u808_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_79a785f7_u0<=1'h0;
else reg_79a785f7_u0<=and_u4087_u0;
end
assign and_u4087_u0=and_u4075_u0&and_u4089_u0;
assign mux_u411_u0=(reg_79a785f7_u0)?mux_u408_u0:syncEnable_u807_u0;
always @(posedge CLK)
begin
if (and_u4089_u0)
syncEnable_u808_u0<=mux_u419_u0;
end
assign and_u4088_u0=and_u4074_u0&and_u4090_u0;
assign mux_u412_u0=(and_delayed_u277_u0)?syncEnable_u809_u0:mux_u410_u0;
assign and_u4089_u0=and_u4073_u0&and_u4090_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u276_u0<=1'h0;
else and_delayed_u276_u0<=and_u4089_u0;
end
always @(posedge CLK)
begin
if (and_u4090_u0)
syncEnable_u809_u0<=mux_u419_u0;
end
assign mux_u413_u0=(and_delayed_u277_u0)?syncEnable_u810_u0:mux_u411_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u277_u0<=1'h0;
else and_delayed_u277_u0<=and_u4088_u0;
end
always @(posedge CLK)
begin
if (and_u4090_u0)
syncEnable_u810_u0<=mux_u418_u0;
end
assign or_u1214_u0=or_u1210_u0|and_u4084_u0;
assign mux_u414_u0=(or_u1210_u0)?1'h1:1'h0;
always @(posedge CLK)
begin
if (block_GO_delayed_u13)
latch_7563f172_reg<=mux_u412_u0;
end
assign latch_7563f172_out=(block_GO_delayed_u13)?mux_u412_u0:latch_7563f172_reg;
assign latch_4c497753_out=(block_GO_delayed_u13)?mux_u413_u0:latch_4c497753_reg;
always @(posedge CLK)
begin
if (block_GO_delayed_u13)
latch_4c497753_reg<=mux_u413_u0;
end
assign mux_u415_u0=(or_u1208_u0)?mux_u405_u0:1'h0;
assign or_u1215_u0=or_u1208_u0|and_u4084_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
block_GO_delayed_u13<=1'h0;
else block_GO_delayed_u13<=and_u4090_u0;
end
assign mux_u416_u0=(or_u1212_u0)?32'h0:add_u575;
assign or_u1216_u0=or_u1212_u0|and_u4082_u0;
assign or_u1217_u0=or_u1209_u0|and_u4084_u0;
assign mux_u417_u0=(or_u1209_u0)?{22'b0, mux_u406_u0[9], 5'b0, mux_u406_u0[3], 3'b0}:32'hffffffff;
assign and_u4090_u0=or_u1218_u0&or_u1218_u0;
assign mux_u418_u0=(loopControl_u10)?fbReg_Out1Portvalue_u5:16'h0;
assign or_u1218_u0=loopControl_u10|reg_4dbfab2c_u0;
assign mux_u419_u0=(loopControl_u10)?fbReg_temp_fsmOldState_resized_LH3_xy_8_u0:32'h0;
always @(posedge CLK)
begin
if (or_u1213_u0)
fbReg_Out1Portvalue_u5<=latch_4c497753_out;
end
always @(posedge CLK)
begin
if (or_u1213_u0)
fbReg_temp_fsmOldState_resized_LH3_xy_8_u0<=latch_7563f172_out;
end
always @(posedge CLK)
begin
if (reg_4dbfab2c_u0)
syncEnable_u811_u0<=RESET;
end
always @(posedge CLK or posedge syncEnable_u811_u0)
begin
if (syncEnable_u811_u0)
loopControl_u10<=1'h0;
else loopControl_u10<=or_u1213_u0;
end
assign mux_u420_u0=(GO)?32'hffffffff:mux_u417_u0;
assign or_u1219_u0=GO|or_u1217_u0;
assign or_u1220_u0=GO|or_u1207_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4dbfab2c_u0<=1'h0;
else reg_4dbfab2c_u0<=reg_585ee52a_u0;
end
assign or_u1221_u0=GO|or_u1216_u0;
assign mux_u421_u0=(GO)?32'h0:mux_u416_u0;
assign mux_u422_u0=(GO)?1'h0:mux_u414_u0;
assign or_u1222_u0=GO|or_u1214_u0;
assign or_u1223_u0=GO|or_u1215_u0;
assign mux_u423_u0=(GO)?1'h0:mux_u415_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_585ee52a_u0<=1'h0;
else reg_585ee52a_u0<=GO;
end
assign RESULT=or_u1220_u0;
assign RESULT_u2370=32'h0;
assign RESULT_u2371=or_u1223_u0;
assign RESULT_u2372=mux_u423_u0;
assign RESULT_u2373=or_u1221_u0;
assign RESULT_u2374=mux_u421_u0;
assign RESULT_u2375=or_u1219_u0;
assign RESULT_u2376=mux_u420_u0;
assign RESULT_u2377=or_u1222_u0;
assign RESULT_u2378=mux_u422_u0;
assign RESULT_u2379=and_u4082_u0;
assign RESULT_u2380=add;
assign RESULT_u2381=3'h1;
assign RESULT_u2382=simplePinWrite_u568;
assign RESULT_u2383=simplePinWrite_u569;
assign RESULT_u2384=simplePinWrite_u570;
assign RESULT_u2385=simplePinWrite;
assign RESULT_u2386=simplePinWrite_u566;
assign RESULT_u2387=simplePinWrite_u567;
assign DONE=1'h0;
endmodule



module resized_LH3_xy_forge_memory_512x16_43(CLK, EN, WE, ADDR, DIN, DOUT, DONE);
input		CLK;
input		EN;
input		WE;
input	[31:0]	ADDR;
input	[15:0]	DIN;
output	[15:0]	DOUT;
output		DONE;
wire		we_0;
wire	[15:0]	pre_dout_0;
wire		we_1;
wire	[15:0]	pre_dout_1;
wire		we_2;
wire	[15:0]	pre_dout_2;
wire		we_3;
wire	[15:0]	pre_dout_3;
reg	[15:0]	mux_out;
reg		wen_done;
assign we_0=WE&(ADDR[31:7]==25'h0);
assign we_1=WE&(ADDR[31:7]==25'h1);
assign we_2=WE&(ADDR[31:7]==25'h2);
assign we_3=WE&(ADDR[31:7]==25'h3);
always @(ADDR or pre_dout_0 or pre_dout_1 or pre_dout_2 or pre_dout_3)
begin
case (ADDR[31:7])25'd0:mux_out=pre_dout_0;
25'd1:mux_out=pre_dout_1;
25'd2:mux_out=pre_dout_2;
25'd3:mux_out=pre_dout_3;
default:mux_out=16'h0;
endcase end
always @(posedge CLK)
begin
wen_done<=WE;
end
assign DOUT=mux_out;
assign DONE=EN&!WE|wen_done;
//  Memory array element: COL: 0, ROW: 0
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_320(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[0]), .O(pre_dout_0[0]));
//  Memory array element: COL: 0, ROW: 1
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_321(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[1]), .O(pre_dout_0[1]));
//  Memory array element: COL: 0, ROW: 2
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_322(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[2]), .O(pre_dout_0[2]));
//  Memory array element: COL: 0, ROW: 3
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_323(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[3]), .O(pre_dout_0[3]));
//  Memory array element: COL: 0, ROW: 4
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_324(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[4]), .O(pre_dout_0[4]));
//  Memory array element: COL: 0, ROW: 5
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_325(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[5]), .O(pre_dout_0[5]));
//  Memory array element: COL: 0, ROW: 6
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_326(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[6]), .O(pre_dout_0[6]));
//  Memory array element: COL: 0, ROW: 7
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_327(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[7]), .O(pre_dout_0[7]));
//  Memory array element: COL: 0, ROW: 8
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_328(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[8]), .O(pre_dout_0[8]));
//  Memory array element: COL: 0, ROW: 9
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_329(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[9]), .O(pre_dout_0[9]));
//  Memory array element: COL: 0, ROW: 10
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_330(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[10]), .O(pre_dout_0[10]));
//  Memory array element: COL: 0, ROW: 11
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_331(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[11]), .O(pre_dout_0[11]));
//  Memory array element: COL: 0, ROW: 12
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_332(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[12]), .O(pre_dout_0[12]));
//  Memory array element: COL: 0, ROW: 13
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_333(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[13]), .O(pre_dout_0[13]));
//  Memory array element: COL: 0, ROW: 14
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_334(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[14]), .O(pre_dout_0[14]));
//  Memory array element: COL: 0, ROW: 15
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_335(.WCLK(CLK), 
  .WE(we_0), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[15]), .O(pre_dout_0[15]));
//  Memory array element: COL: 1, ROW: 0
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_336(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[0]), .O(pre_dout_1[0]));
//  Memory array element: COL: 1, ROW: 1
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_337(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[1]), .O(pre_dout_1[1]));
//  Memory array element: COL: 1, ROW: 2
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_338(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[2]), .O(pre_dout_1[2]));
//  Memory array element: COL: 1, ROW: 3
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_339(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[3]), .O(pre_dout_1[3]));
//  Memory array element: COL: 1, ROW: 4
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_340(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[4]), .O(pre_dout_1[4]));
//  Memory array element: COL: 1, ROW: 5
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_341(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[5]), .O(pre_dout_1[5]));
//  Memory array element: COL: 1, ROW: 6
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_342(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[6]), .O(pre_dout_1[6]));
//  Memory array element: COL: 1, ROW: 7
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_343(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[7]), .O(pre_dout_1[7]));
//  Memory array element: COL: 1, ROW: 8
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_344(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[8]), .O(pre_dout_1[8]));
//  Memory array element: COL: 1, ROW: 9
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_345(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[9]), .O(pre_dout_1[9]));
//  Memory array element: COL: 1, ROW: 10
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_346(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[10]), .O(pre_dout_1[10]));
//  Memory array element: COL: 1, ROW: 11
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_347(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[11]), .O(pre_dout_1[11]));
//  Memory array element: COL: 1, ROW: 12
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_348(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[12]), .O(pre_dout_1[12]));
//  Memory array element: COL: 1, ROW: 13
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_349(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[13]), .O(pre_dout_1[13]));
//  Memory array element: COL: 1, ROW: 14
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_350(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[14]), .O(pre_dout_1[14]));
//  Memory array element: COL: 1, ROW: 15
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_351(.WCLK(CLK), 
  .WE(we_1), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[15]), .O(pre_dout_1[15]));
//  Memory array element: COL: 2, ROW: 0
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_352(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[0]), .O(pre_dout_2[0]));
//  Memory array element: COL: 2, ROW: 1
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_353(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[1]), .O(pre_dout_2[1]));
//  Memory array element: COL: 2, ROW: 2
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_354(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[2]), .O(pre_dout_2[2]));
//  Memory array element: COL: 2, ROW: 3
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_355(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[3]), .O(pre_dout_2[3]));
//  Memory array element: COL: 2, ROW: 4
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_356(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[4]), .O(pre_dout_2[4]));
//  Memory array element: COL: 2, ROW: 5
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_357(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[5]), .O(pre_dout_2[5]));
//  Memory array element: COL: 2, ROW: 6
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_358(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[6]), .O(pre_dout_2[6]));
//  Memory array element: COL: 2, ROW: 7
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_359(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[7]), .O(pre_dout_2[7]));
//  Memory array element: COL: 2, ROW: 8
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_360(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[8]), .O(pre_dout_2[8]));
//  Memory array element: COL: 2, ROW: 9
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_361(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[9]), .O(pre_dout_2[9]));
//  Memory array element: COL: 2, ROW: 10
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_362(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[10]), .O(pre_dout_2[10]));
//  Memory array element: COL: 2, ROW: 11
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_363(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[11]), .O(pre_dout_2[11]));
//  Memory array element: COL: 2, ROW: 12
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_364(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[12]), .O(pre_dout_2[12]));
//  Memory array element: COL: 2, ROW: 13
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_365(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[13]), .O(pre_dout_2[13]));
//  Memory array element: COL: 2, ROW: 14
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_366(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[14]), .O(pre_dout_2[14]));
//  Memory array element: COL: 2, ROW: 15
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_367(.WCLK(CLK), 
  .WE(we_2), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[15]), .O(pre_dout_2[15]));
//  Memory array element: COL: 3, ROW: 0
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_368(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[0]), .O(pre_dout_3[0]));
//  Memory array element: COL: 3, ROW: 1
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_369(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[1]), .O(pre_dout_3[1]));
//  Memory array element: COL: 3, ROW: 2
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_370(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[2]), .O(pre_dout_3[2]));
//  Memory array element: COL: 3, ROW: 3
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_371(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[3]), .O(pre_dout_3[3]));
//  Memory array element: COL: 3, ROW: 4
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_372(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[4]), .O(pre_dout_3[4]));
//  Memory array element: COL: 3, ROW: 5
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_373(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[5]), .O(pre_dout_3[5]));
//  Memory array element: COL: 3, ROW: 6
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_374(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[6]), .O(pre_dout_3[6]));
//  Memory array element: COL: 3, ROW: 7
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_375(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[7]), .O(pre_dout_3[7]));
//  Memory array element: COL: 3, ROW: 8
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_376(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[8]), .O(pre_dout_3[8]));
//  Memory array element: COL: 3, ROW: 9
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_377(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[9]), .O(pre_dout_3[9]));
//  Memory array element: COL: 3, ROW: 10
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_378(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[10]), .O(pre_dout_3[10]));
//  Memory array element: COL: 3, ROW: 11
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_379(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[11]), .O(pre_dout_3[11]));
//  Memory array element: COL: 3, ROW: 12
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_380(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[12]), .O(pre_dout_3[12]));
//  Memory array element: COL: 3, ROW: 13
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_381(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[13]), .O(pre_dout_3[13]));
//  Memory array element: COL: 3, ROW: 14
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_382(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[14]), .O(pre_dout_3[14]));
//  Memory array element: COL: 3, ROW: 15
//  Initialization of LUT ram is accomplished through explicit parameter
// setting.
RAM128X1S#(.INIT(128'h00000000000000000000000000000000))RAM128X1S_instance_383(.WCLK(CLK), 
  .WE(we_3), .A0(ADDR[0]), .A1(ADDR[1]), .A2(ADDR[2]), .A3(ADDR[3]), .A4(ADDR[4]), .A5(ADDR[5]), 
  .A6(ADDR[6]), .D(DIN[15]), .O(pre_dout_3[15]));
endmodule



module resized_LH3_xy_structuralmemory_5a4854c1_(CLK_u23, bus_4424cad2_, bus_287c41c7_, bus_66538fba_, bus_793de9c2_, bus_1f47f383_, bus_462ad95f_, bus_6f4f27ab_, bus_5cd62f8e_);
input		CLK_u23;
input		bus_4424cad2_;
input	[31:0]	bus_287c41c7_;
input	[2:0]	bus_66538fba_;
input		bus_793de9c2_;
input		bus_1f47f383_;
input	[15:0]	bus_462ad95f_;
output	[15:0]	bus_6f4f27ab_;
output		bus_5cd62f8e_;
wire		or_34c2bb42_u0;
reg		logicalMem_7d94c52d_we_delay0_u0=1'h0;
wire		or_5b9ccd5e_u0;
wire		not_7a2fbd81_u0;
wire	[15:0]	bus_5f7afa32_;
wire		and_2a77a863_u0;
assign or_34c2bb42_u0=bus_793de9c2_|bus_1f47f383_;
always @(posedge CLK_u23 or posedge bus_4424cad2_)
begin
if (bus_4424cad2_)
logicalMem_7d94c52d_we_delay0_u0<=1'h0;
else logicalMem_7d94c52d_we_delay0_u0<=bus_1f47f383_;
end
assign or_5b9ccd5e_u0=and_2a77a863_u0|logicalMem_7d94c52d_we_delay0_u0;
assign not_7a2fbd81_u0=~bus_1f47f383_;
assign bus_6f4f27ab_=bus_5f7afa32_;
assign bus_5cd62f8e_=or_5b9ccd5e_u0;
resized_LH3_xy_forge_memory_512x16_43 resized_LH3_xy_forge_memory_512x16_43_instance0(.CLK(CLK_u23), 
  .EN(or_34c2bb42_u0), .WE(bus_1f47f383_), .ADDR(bus_287c41c7_), .DIN(bus_462ad95f_), 
  .DOUT(bus_5f7afa32_), .DONE());
assign and_2a77a863_u0=bus_793de9c2_&not_7a2fbd81_u0;
endmodule



module resized_LH3_xy_simplememoryreferee_4dbf2a2f_(bus_170ffe51_, bus_2bdc80e5_, bus_5068a6cf_, bus_4a24c1e1_, bus_71489945_, bus_0668b190_, bus_69dc047c_, bus_419996e9_, bus_309461d8_, bus_0943531d_, bus_1bce23d3_, bus_6d8c43ff_, bus_67ef8aa5_, bus_3032e61d_, bus_7a45fad8_, bus_7927363a_, bus_1598a4d3_, bus_39892bbf_, bus_604acdab_, bus_1310b3e4_, bus_4497015b_, bus_5d365df5_, bus_0859aa58_, bus_4eb99653_);
input		bus_170ffe51_;
input		bus_2bdc80e5_;
input		bus_5068a6cf_;
input	[15:0]	bus_4a24c1e1_;
input		bus_71489945_;
input	[15:0]	bus_0668b190_;
input	[31:0]	bus_69dc047c_;
input	[2:0]	bus_419996e9_;
input		bus_309461d8_;
input	[15:0]	bus_0943531d_;
input	[31:0]	bus_1bce23d3_;
input	[2:0]	bus_6d8c43ff_;
input		bus_67ef8aa5_;
input	[31:0]	bus_3032e61d_;
input	[2:0]	bus_7a45fad8_;
output	[15:0]	bus_7927363a_;
output	[31:0]	bus_1598a4d3_;
output		bus_39892bbf_;
output		bus_604acdab_;
output	[2:0]	bus_1310b3e4_;
output		bus_4497015b_;
output		bus_5d365df5_;
output	[15:0]	bus_0859aa58_;
output		bus_4eb99653_;
wire		or_4bd6c336_u0;
reg		done_qual_u225=1'h0;
wire		and_0fde70f5_u0;
wire	[15:0]	mux_78783254_u0;
reg		done_qual_u226_u0=1'h0;
wire		not_2ac81507_u0;
wire		or_3daf991f_u0;
wire		and_2cf2f682_u0;
wire		and_23a71716_u0;
wire		or_62da7629_u0;
wire		not_0fa24836_u0;
wire		not_5623a675_u0;
wire		or_6356b4ce_u0;
wire	[31:0]	mux_54fcb425_u0;
wire		or_72099774_u0;
reg		done_qual_u227_u0=1'h0;
assign or_4bd6c336_u0=bus_67ef8aa5_|done_qual_u225;
always @(posedge bus_170ffe51_)
begin
if (bus_2bdc80e5_)
done_qual_u225<=1'h0;
else done_qual_u225<=bus_67ef8aa5_;
end
assign and_0fde70f5_u0=or_4bd6c336_u0&bus_5068a6cf_;
assign mux_78783254_u0=(bus_71489945_)?bus_0668b190_:bus_0943531d_;
assign bus_7927363a_=mux_78783254_u0;
assign bus_1598a4d3_=mux_54fcb425_u0;
assign bus_39892bbf_=or_72099774_u0;
assign bus_604acdab_=or_62da7629_u0;
assign bus_1310b3e4_=3'h1;
assign bus_4497015b_=and_23a71716_u0;
assign bus_5d365df5_=and_2cf2f682_u0;
assign bus_0859aa58_=bus_4a24c1e1_;
assign bus_4eb99653_=and_0fde70f5_u0;
always @(posedge bus_170ffe51_)
begin
if (bus_2bdc80e5_)
done_qual_u226_u0<=1'h0;
else done_qual_u226_u0<=bus_309461d8_;
end
assign not_2ac81507_u0=~bus_5068a6cf_;
assign or_3daf991f_u0=bus_71489945_|done_qual_u227_u0;
assign and_2cf2f682_u0=or_6356b4ce_u0&bus_5068a6cf_;
assign and_23a71716_u0=or_3daf991f_u0&bus_5068a6cf_;
assign or_62da7629_u0=bus_71489945_|bus_309461d8_|bus_67ef8aa5_;
assign not_0fa24836_u0=~bus_5068a6cf_;
assign not_5623a675_u0=~bus_5068a6cf_;
assign or_6356b4ce_u0=bus_309461d8_|done_qual_u226_u0;
assign mux_54fcb425_u0=({32{bus_71489945_}}&bus_69dc047c_)|({32{bus_309461d8_}}&bus_1bce23d3_)|({32{bus_67ef8aa5_}}&bus_3032e61d_);
assign or_72099774_u0=bus_71489945_|bus_309461d8_;
always @(posedge bus_170ffe51_)
begin
if (bus_2bdc80e5_)
done_qual_u227_u0<=1'h0;
else done_qual_u227_u0<=bus_71489945_;
end
endmodule



module resized_LH3_xy_globalreset_physical_6b469655_(bus_7bfcb29f_, bus_21c9004a_, bus_45a18503_);
input		bus_7bfcb29f_;
input		bus_21c9004a_;
output		bus_45a18503_;
reg		cross_u43=1'h0;
reg		glitch_u43=1'h0;
reg		sample_u43=1'h0;
wire		not_0124b7cf_u0;
wire		and_7f4d6041_u0;
wire		or_0b0d2041_u0;
reg		final_u43=1'h1;
always @(posedge bus_7bfcb29f_)
begin
cross_u43<=sample_u43;
end
always @(posedge bus_7bfcb29f_)
begin
glitch_u43<=cross_u43;
end
always @(posedge bus_7bfcb29f_)
begin
sample_u43<=1'h1;
end
assign not_0124b7cf_u0=~and_7f4d6041_u0;
assign and_7f4d6041_u0=cross_u43&glitch_u43;
assign or_0b0d2041_u0=bus_21c9004a_|final_u43;
assign bus_45a18503_=or_0b0d2041_u0;
always @(posedge bus_7bfcb29f_)
begin
final_u43<=not_0124b7cf_u0;
end
endmodule



module resized_LH3_xy_Kicker_47(CLK, RESET, bus_3606f0fa_);
input		CLK;
input		RESET;
output		bus_3606f0fa_;
reg		kicker_res=1'h0;
wire		bus_352dd25f_;
wire		bus_185364c5_;
reg		kicker_1=1'h0;
reg		kicker_2=1'h0;
wire		bus_4774a6ff_;
wire		bus_45aca703_;
assign bus_3606f0fa_=kicker_res;
always @(posedge CLK)
begin
kicker_res<=bus_4774a6ff_;
end
assign bus_352dd25f_=~RESET;
assign bus_185364c5_=bus_352dd25f_&kicker_1;
always @(posedge CLK)
begin
kicker_1<=bus_352dd25f_;
end
always @(posedge CLK)
begin
kicker_2<=bus_185364c5_;
end
assign bus_4774a6ff_=kicker_1&bus_352dd25f_&bus_45aca703_;
assign bus_45aca703_=~kicker_2;
endmodule



module resized_LH3_xy_endianswapper_5dd691e5_(endianswapper_5dd691e5_in, endianswapper_5dd691e5_out);
input	[15:0]	endianswapper_5dd691e5_in;
output	[15:0]	endianswapper_5dd691e5_out;
assign endianswapper_5dd691e5_out=endianswapper_5dd691e5_in;
endmodule



module resized_LH3_xy_endianswapper_3372e3cb_(endianswapper_3372e3cb_in, endianswapper_3372e3cb_out);
input	[15:0]	endianswapper_3372e3cb_in;
output	[15:0]	endianswapper_3372e3cb_out;
assign endianswapper_3372e3cb_out=endianswapper_3372e3cb_in;
endmodule



module resized_LH3_xy_stateVar_x(bus_21f26c1b_, bus_27078042_, bus_318dd820_, bus_18336d09_, bus_26bd9abe_, bus_49e109b4_, bus_33af6980_);
input		bus_21f26c1b_;
input		bus_27078042_;
input		bus_318dd820_;
input	[15:0]	bus_18336d09_;
input		bus_26bd9abe_;
input	[15:0]	bus_49e109b4_;
output	[15:0]	bus_33af6980_;
wire	[15:0]	endianswapper_5dd691e5_out;
reg	[15:0]	stateVar_x_u5=16'h0;
wire		or_4138bc00_u0;
wire	[15:0]	endianswapper_3372e3cb_out;
wire	[15:0]	mux_4635dc2e_u0;
resized_LH3_xy_endianswapper_5dd691e5_ resized_LH3_xy_endianswapper_5dd691e5__1(.endianswapper_5dd691e5_in(mux_4635dc2e_u0), 
  .endianswapper_5dd691e5_out(endianswapper_5dd691e5_out));
assign bus_33af6980_=endianswapper_3372e3cb_out;
always @(posedge bus_21f26c1b_ or posedge bus_27078042_)
begin
if (bus_27078042_)
stateVar_x_u5<=16'h0;
else if (or_4138bc00_u0)
stateVar_x_u5<=endianswapper_5dd691e5_out;
end
assign or_4138bc00_u0=bus_318dd820_|bus_26bd9abe_;
resized_LH3_xy_endianswapper_3372e3cb_ resized_LH3_xy_endianswapper_3372e3cb__1(.endianswapper_3372e3cb_in(stateVar_x_u5), 
  .endianswapper_3372e3cb_out(endianswapper_3372e3cb_out));
assign mux_4635dc2e_u0=(bus_318dd820_)?bus_18336d09_:16'h0;
endmodule



module resized_LH3_xy_endianswapper_30af27d9_(endianswapper_30af27d9_in, endianswapper_30af27d9_out);
input	[15:0]	endianswapper_30af27d9_in;
output	[15:0]	endianswapper_30af27d9_out;
assign endianswapper_30af27d9_out=endianswapper_30af27d9_in;
endmodule



module resized_LH3_xy_endianswapper_049793d8_(endianswapper_049793d8_in, endianswapper_049793d8_out);
input	[15:0]	endianswapper_049793d8_in;
output	[15:0]	endianswapper_049793d8_out;
assign endianswapper_049793d8_out=endianswapper_049793d8_in;
endmodule



module resized_LH3_xy_stateVar_rowRepeated(bus_45f031f5_, bus_1b617bad_, bus_3bba85fa_, bus_6fadc4af_, bus_4ba53be4_, bus_3e7ecbe0_, bus_5e36be26_);
input		bus_45f031f5_;
input		bus_1b617bad_;
input		bus_3bba85fa_;
input	[15:0]	bus_6fadc4af_;
input		bus_4ba53be4_;
input	[15:0]	bus_3e7ecbe0_;
output	[15:0]	bus_5e36be26_;
wire		or_6d238117_u0;
reg	[15:0]	stateVar_rowRepeated_u5=16'h1;
wire	[15:0]	endianswapper_30af27d9_out;
wire	[15:0]	mux_5b98ae35_u0;
wire	[15:0]	endianswapper_049793d8_out;
assign bus_5e36be26_=endianswapper_30af27d9_out;
assign or_6d238117_u0=bus_3bba85fa_|bus_4ba53be4_;
always @(posedge bus_45f031f5_ or posedge bus_1b617bad_)
begin
if (bus_1b617bad_)
stateVar_rowRepeated_u5<=16'h1;
else if (or_6d238117_u0)
stateVar_rowRepeated_u5<=endianswapper_049793d8_out;
end
resized_LH3_xy_endianswapper_30af27d9_ resized_LH3_xy_endianswapper_30af27d9__1(.endianswapper_30af27d9_in(stateVar_rowRepeated_u5), 
  .endianswapper_30af27d9_out(endianswapper_30af27d9_out));
assign mux_5b98ae35_u0=(bus_3bba85fa_)?bus_6fadc4af_:16'h1;
resized_LH3_xy_endianswapper_049793d8_ resized_LH3_xy_endianswapper_049793d8__1(.endianswapper_049793d8_in(mux_5b98ae35_u0), 
  .endianswapper_049793d8_out(endianswapper_049793d8_out));
endmodule



module resized_LH3_xy_endianswapper_04967a21_(endianswapper_04967a21_in, endianswapper_04967a21_out);
input	[31:0]	endianswapper_04967a21_in;
output	[31:0]	endianswapper_04967a21_out;
assign endianswapper_04967a21_out=32'h0;
endmodule



module resized_LH3_xy_endianswapper_4dbbaf73_(endianswapper_4dbbaf73_in, endianswapper_4dbbaf73_out);
input	[31:0]	endianswapper_4dbbaf73_in;
output	[31:0]	endianswapper_4dbbaf73_out;
assign endianswapper_4dbbaf73_out=32'h0;
endmodule



module resized_LH3_xy_stateVar_fsmOldState_resized_LH3_xy(bus_1e850958_, bus_0fe2bf8a_, bus_2d9446c1_, bus_0169b7ea_, bus_48c16de3_);
input		bus_1e850958_;
input		bus_0fe2bf8a_;
input		bus_2d9446c1_;
input	[31:0]	bus_0169b7ea_;
output	[31:0]	bus_48c16de3_;
wire	[31:0]	endianswapper_04967a21_out;
wire	[31:0]	endianswapper_4dbbaf73_out;
assign bus_48c16de3_=32'h0;
resized_LH3_xy_endianswapper_04967a21_ resized_LH3_xy_endianswapper_04967a21__1(.endianswapper_04967a21_in(32'h0), 
  .endianswapper_04967a21_out(endianswapper_04967a21_out));
resized_LH3_xy_endianswapper_4dbbaf73_ resized_LH3_xy_endianswapper_4dbbaf73__1(.endianswapper_4dbbaf73_in(32'h0), 
  .endianswapper_4dbbaf73_out(endianswapper_4dbbaf73_out));
endmodule



module resized_LH3_xy_simplememoryreferee_10f2e65e_(bus_095cf1de_, bus_1d16e5f4_, bus_15440525_, bus_1f52af7b_, bus_5d57546f_, bus_23881311_, bus_385fd4fe_, bus_074a4e9c_, bus_0109f5e5_, bus_38ee4680_, bus_55728af0_, bus_07b29725_, bus_36c9b0d0_, bus_2f725b02_, bus_30f6e3b0_, bus_6620e554_, bus_38031f96_, bus_21d6a5fd_, bus_12a86ec5_);
input		bus_095cf1de_;
input		bus_1d16e5f4_;
input		bus_15440525_;
input	[15:0]	bus_1f52af7b_;
input		bus_5d57546f_;
input	[15:0]	bus_23881311_;
input	[31:0]	bus_385fd4fe_;
input	[2:0]	bus_074a4e9c_;
input		bus_0109f5e5_;
input	[31:0]	bus_38ee4680_;
input	[2:0]	bus_55728af0_;
output	[15:0]	bus_07b29725_;
output	[31:0]	bus_36c9b0d0_;
output		bus_2f725b02_;
output		bus_30f6e3b0_;
output	[2:0]	bus_6620e554_;
output		bus_38031f96_;
output	[15:0]	bus_21d6a5fd_;
output		bus_12a86ec5_;
wire	[15:0]	mux_6b21cce1_u0;
reg		done_qual_u228_u0=1'h0;
wire		not_5ab00bf8_u0;
wire		and_2d5f16d4_u0;
wire	[31:0]	mux_5e0ce61c_u0;
wire		not_4a89cbb8_u0;
wire		or_41fd252e_u0;
wire		or_6b43631a_u0;
wire		or_5f6046bb_u0;
wire		and_78a1563c_u0;
reg		done_qual_u229_u0=1'h0;
assign mux_6b21cce1_u0=({16{bus_5d57546f_}}&bus_23881311_);
always @(posedge bus_095cf1de_)
begin
if (bus_1d16e5f4_)
done_qual_u228_u0<=1'h0;
else done_qual_u228_u0<=bus_0109f5e5_;
end
assign not_5ab00bf8_u0=~bus_15440525_;
assign and_2d5f16d4_u0=or_5f6046bb_u0&bus_15440525_;
assign mux_5e0ce61c_u0=(bus_5d57546f_)?bus_385fd4fe_:bus_38ee4680_;
assign not_4a89cbb8_u0=~bus_15440525_;
assign or_41fd252e_u0=bus_0109f5e5_|done_qual_u228_u0;
assign or_6b43631a_u0=bus_5d57546f_|bus_0109f5e5_;
assign or_5f6046bb_u0=bus_5d57546f_|done_qual_u229_u0;
assign bus_07b29725_=mux_6b21cce1_u0;
assign bus_36c9b0d0_=mux_5e0ce61c_u0;
assign bus_2f725b02_=bus_5d57546f_;
assign bus_30f6e3b0_=or_6b43631a_u0;
assign bus_6620e554_=3'h1;
assign bus_38031f96_=and_2d5f16d4_u0;
assign bus_21d6a5fd_=bus_1f52af7b_;
assign bus_12a86ec5_=and_78a1563c_u0;
assign and_78a1563c_u0=or_41fd252e_u0&bus_15440525_;
always @(posedge bus_095cf1de_)
begin
if (bus_1d16e5f4_)
done_qual_u229_u0<=1'h0;
else done_qual_u229_u0<=bus_5d57546f_;
end
endmodule



module resized_LH3_xy_endianswapper_28a15479_(endianswapper_28a15479_in, endianswapper_28a15479_out);
input		endianswapper_28a15479_in;
output		endianswapper_28a15479_out;
assign endianswapper_28a15479_out=endianswapper_28a15479_in;
endmodule



module resized_LH3_xy_endianswapper_0b3c9987_(endianswapper_0b3c9987_in, endianswapper_0b3c9987_out);
input		endianswapper_0b3c9987_in;
output		endianswapper_0b3c9987_out;
assign endianswapper_0b3c9987_out=endianswapper_0b3c9987_in;
endmodule



module resized_LH3_xy_stateVar_fsmState_resized_LH3_xy(bus_35a4b222_, bus_1fa30b0d_, bus_7894e09d_, bus_6f4dfd67_, bus_61fe06bb_);
input		bus_35a4b222_;
input		bus_1fa30b0d_;
input		bus_7894e09d_;
input		bus_6f4dfd67_;
output		bus_61fe06bb_;
wire		endianswapper_28a15479_out;
reg		stateVar_fsmState_resized_LH3_xy_u0=1'h0;
wire		endianswapper_0b3c9987_out;
resized_LH3_xy_endianswapper_28a15479_ resized_LH3_xy_endianswapper_28a15479__1(.endianswapper_28a15479_in(bus_6f4dfd67_), 
  .endianswapper_28a15479_out(endianswapper_28a15479_out));
always @(posedge bus_35a4b222_ or posedge bus_1fa30b0d_)
begin
if (bus_1fa30b0d_)
stateVar_fsmState_resized_LH3_xy_u0<=1'h0;
else if (bus_7894e09d_)
stateVar_fsmState_resized_LH3_xy_u0<=endianswapper_28a15479_out;
end
resized_LH3_xy_endianswapper_0b3c9987_ resized_LH3_xy_endianswapper_0b3c9987__1(.endianswapper_0b3c9987_in(stateVar_fsmState_resized_LH3_xy_u0), 
  .endianswapper_0b3c9987_out(endianswapper_0b3c9987_out));
assign bus_61fe06bb_=endianswapper_0b3c9987_out;
endmodule



module resized_LH3_xy_repeatRowExpanded(CLK, RESET, GO, port_7ef0238d_, port_138273d0_, port_183b6d71_, port_466e1c3e_, RESULT, RESULT_u2388, RESULT_u2389, RESULT_u2390, RESULT_u2391, RESULT_u2392, RESULT_u2393, RESULT_u2394, RESULT_u2395, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_7ef0238d_;
input		port_138273d0_;
input		port_183b6d71_;
input	[15:0]	port_466e1c3e_;
output		RESULT;
output	[15:0]	RESULT_u2388;
output		RESULT_u2389;
output	[31:0]	RESULT_u2390;
output	[15:0]	RESULT_u2391;
output	[2:0]	RESULT_u2392;
output		RESULT_u2393;
output	[31:0]	RESULT_u2394;
output	[2:0]	RESULT_u2395;
output		DONE;
wire	[15:0]	add;
wire	[31:0]	add_u576;
wire		and_u4091_u0;
wire	[31:0]	add_u577;
wire		or_u1224_u0;
reg		reg_080c828b_u0=1'h0;
wire		and_u4092_u0;
wire	[31:0]	add_u578;
reg	[31:0]	syncEnable_u812=32'h0;
wire		and_u4093_u0;
wire		lessThan;
wire signed	[31:0]	lessThan_b_signed;
wire signed	[31:0]	lessThan_a_signed;
wire		not_u653_u0;
wire		and_u4094_u0;
wire		and_u4095_u0;
reg		and_delayed_u278=1'h0;
wire		and_u4096_u0;
wire	[31:0]	mux_u424;
wire		or_u1225_u0;
reg		reg_6e40ff8d_u0=1'h0;
assign add=port_7ef0238d_+16'h1;
assign add_u576=mux_u424+32'h0;
assign and_u4091_u0=and_u4093_u0&port_183b6d71_;
assign add_u577=mux_u424+32'h0;
assign or_u1224_u0=and_u4092_u0|RESET;
always @(posedge CLK or posedge and_u4093_u0 or posedge or_u1224_u0)
begin
if (or_u1224_u0)
reg_080c828b_u0<=1'h0;
else if (and_u4093_u0)
reg_080c828b_u0<=1'h1;
else reg_080c828b_u0<=reg_080c828b_u0;
end
assign and_u4092_u0=reg_080c828b_u0&port_138273d0_;
assign add_u578=mux_u424+32'h1;
always @(posedge CLK)
begin
if (and_u4093_u0)
syncEnable_u812<=add_u578;
end
assign and_u4093_u0=and_u4094_u0&or_u1225_u0;
assign lessThan_a_signed=mux_u424;
assign lessThan_b_signed=32'h200;
assign lessThan=lessThan_a_signed<lessThan_b_signed;
assign not_u653_u0=~lessThan;
assign and_u4094_u0=or_u1225_u0&lessThan;
assign and_u4095_u0=or_u1225_u0&not_u653_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u278<=1'h0;
else and_delayed_u278<=and_u4093_u0;
end
assign and_u4096_u0=and_u4095_u0&or_u1225_u0;
assign mux_u424=(and_delayed_u278)?syncEnable_u812:32'h0;
assign or_u1225_u0=and_delayed_u278|reg_6e40ff8d_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_6e40ff8d_u0<=1'h0;
else reg_6e40ff8d_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u2388=add;
assign RESULT_u2389=and_u4093_u0;
assign RESULT_u2390=add_u577;
assign RESULT_u2391=port_466e1c3e_;
assign RESULT_u2392=3'h1;
assign RESULT_u2393=and_u4093_u0;
assign RESULT_u2394=add_u576;
assign RESULT_u2395=3'h1;
assign DONE=and_u4096_u0;
endmodule



module resized_LH3_xy_endianswapper_3295ad84_(endianswapper_3295ad84_in, endianswapper_3295ad84_out);
input	[31:0]	endianswapper_3295ad84_in;
output	[31:0]	endianswapper_3295ad84_out;
assign endianswapper_3295ad84_out=endianswapper_3295ad84_in;
endmodule



module resized_LH3_xy_endianswapper_6da49600_(endianswapper_6da49600_in, endianswapper_6da49600_out);
input	[31:0]	endianswapper_6da49600_in;
output	[31:0]	endianswapper_6da49600_out;
assign endianswapper_6da49600_out=endianswapper_6da49600_in;
endmodule



module resized_LH3_xy_stateVar_Out1TokenIndex(bus_240b7571_, bus_2effa3d4_, bus_69e423e6_, bus_45898356_, bus_32281ea7_);
input		bus_240b7571_;
input		bus_2effa3d4_;
input		bus_69e423e6_;
input	[31:0]	bus_45898356_;
output	[31:0]	bus_32281ea7_;
wire	[31:0]	endianswapper_3295ad84_out;
reg	[31:0]	stateVar_Out1TokenIndex_u5=32'h0;
wire	[31:0]	endianswapper_6da49600_out;
resized_LH3_xy_endianswapper_3295ad84_ resized_LH3_xy_endianswapper_3295ad84__1(.endianswapper_3295ad84_in(bus_45898356_), 
  .endianswapper_3295ad84_out(endianswapper_3295ad84_out));
always @(posedge bus_240b7571_ or posedge bus_2effa3d4_)
begin
if (bus_2effa3d4_)
stateVar_Out1TokenIndex_u5<=32'h0;
else if (bus_69e423e6_)
stateVar_Out1TokenIndex_u5<=endianswapper_3295ad84_out;
end
resized_LH3_xy_endianswapper_6da49600_ resized_LH3_xy_endianswapper_6da49600__1(.endianswapper_6da49600_in(stateVar_Out1TokenIndex_u5), 
  .endianswapper_6da49600_out(endianswapper_6da49600_out));
assign bus_32281ea7_=endianswapper_6da49600_out;
endmodule



module resized_LH3_xy_reset(CLK, RESET, GO, RESULT, RESULT_u2396, RESULT_u2397, RESULT_u2398, DONE);
input		CLK;
input		RESET;
input		GO;
output		RESULT;
output	[15:0]	RESULT_u2396;
output		RESULT_u2397;
output	[15:0]	RESULT_u2398;
output		DONE;
reg		reg_453f5f2b_u0=1'h0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_453f5f2b_u0<=1'h0;
else reg_453f5f2b_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u2396=16'h1;
assign RESULT_u2397=GO;
assign RESULT_u2398=16'h0;
assign DONE=reg_453f5f2b_u0;
endmodule



module resized_LH3_xy_endianswapper_65eb4a7b_(endianswapper_65eb4a7b_in, endianswapper_65eb4a7b_out);
input	[31:0]	endianswapper_65eb4a7b_in;
output	[31:0]	endianswapper_65eb4a7b_out;
assign endianswapper_65eb4a7b_out=endianswapper_65eb4a7b_in;
endmodule



module resized_LH3_xy_endianswapper_4182fed0_(endianswapper_4182fed0_in, endianswapper_4182fed0_out);
input	[31:0]	endianswapper_4182fed0_in;
output	[31:0]	endianswapper_4182fed0_out;
assign endianswapper_4182fed0_out=endianswapper_4182fed0_in;
endmodule



module resized_LH3_xy_stateVar_Out1MaxTokenIndex(bus_7dd8451b_, bus_6e8b3703_, bus_185d6703_, bus_10961150_, bus_14dbd04d_);
input		bus_7dd8451b_;
input		bus_6e8b3703_;
input		bus_185d6703_;
input	[31:0]	bus_10961150_;
output	[31:0]	bus_14dbd04d_;
wire	[31:0]	endianswapper_65eb4a7b_out;
reg	[31:0]	stateVar_Out1MaxTokenIndex_u5=32'h0;
wire	[31:0]	endianswapper_4182fed0_out;
resized_LH3_xy_endianswapper_65eb4a7b_ resized_LH3_xy_endianswapper_65eb4a7b__1(.endianswapper_65eb4a7b_in(stateVar_Out1MaxTokenIndex_u5), 
  .endianswapper_65eb4a7b_out(endianswapper_65eb4a7b_out));
always @(posedge bus_7dd8451b_ or posedge bus_6e8b3703_)
begin
if (bus_6e8b3703_)
stateVar_Out1MaxTokenIndex_u5<=32'h0;
else if (bus_185d6703_)
stateVar_Out1MaxTokenIndex_u5<=endianswapper_4182fed0_out;
end
resized_LH3_xy_endianswapper_4182fed0_ resized_LH3_xy_endianswapper_4182fed0__1(.endianswapper_4182fed0_in(bus_10961150_), 
  .endianswapper_4182fed0_out(endianswapper_4182fed0_out));
assign bus_14dbd04d_=endianswapper_65eb4a7b_out;
endmodule



module resized_LH3_xy_stateVar_Out1PortEnable(bus_66c9187f_, bus_7bb89c8a_, bus_016a15f2_, bus_10ad7aff_, bus_07319e33_);
input		bus_66c9187f_;
input		bus_7bb89c8a_;
input		bus_016a15f2_;
input		bus_10ad7aff_;
output		bus_07319e33_;
reg		stateVar_Out1PortEnable_u5=1'h0;
assign bus_07319e33_=stateVar_Out1PortEnable_u5;
always @(posedge bus_66c9187f_ or posedge bus_7bb89c8a_)
begin
if (bus_7bb89c8a_)
stateVar_Out1PortEnable_u5<=1'h0;
else if (bus_016a15f2_)
stateVar_Out1PortEnable_u5<=bus_10ad7aff_;
end
endmodule



module resized_LH3_xy_consumeRow(CLK, RESET, GO, port_7ee25a17_, port_00eaa84f_, port_4bf12c4e_, port_0266fa2c_, RESULT, RESULT_u2399, RESULT_u2400, RESULT_u2401, RESULT_u2402, RESULT_u2403, RESULT_u2404, RESULT_u2405, RESULT_u2406, RESULT_u2407, RESULT_u2408, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_7ee25a17_;
input		port_00eaa84f_;
input		port_4bf12c4e_;
input	[15:0]	port_0266fa2c_;
output		RESULT;
output	[15:0]	RESULT_u2399;
output		RESULT_u2400;
output	[31:0]	RESULT_u2401;
output	[15:0]	RESULT_u2402;
output	[2:0]	RESULT_u2403;
output		RESULT_u2404;
output	[31:0]	RESULT_u2405;
output	[15:0]	RESULT_u2406;
output	[2:0]	RESULT_u2407;
output		RESULT_u2408;
output		DONE;
wire		simplePinWrite;
wire signed	[16:0]	lessThanEqualTo_a_signed;
wire		lessThanEqualTo;
wire signed	[16:0]	lessThanEqualTo_b_signed;
wire		and_u4097_u0;
wire		not_u654_u0;
wire		and_u4098_u0;
reg		reg_4a35a071_u0=1'h0;
wire		and_u4099_u0;
wire		and_u4100_u0;
wire	[31:0]	add;
wire	[31:0]	add_u579;
reg		reg_6d0dbf08_u0=1'h0;
wire		and_u4101_u0;
wire		or_u1226_u0;
wire	[15:0]	add_u580;
reg	[15:0]	syncEnable_u813=16'h0;
wire	[15:0]	mux_u425;
wire		or_u1227_u0;
wire	[15:0]	latch_43b8c804_out;
reg	[15:0]	latch_43b8c804_reg=16'h0;
wire	[15:0]	add_u581;
wire		and_u4102_u0;
wire signed	[16:0]	lessThanEqualTo_u5_a_signed;
wire signed	[16:0]	lessThanEqualTo_u5_b_signed;
wire		lessThanEqualTo_u5;
wire		and_u4103_u0;
wire		not_u655_u0;
wire		and_u4104_u0;
reg		and_delayed_u279=1'h0;
wire	[15:0]	subtract;
wire	[31:0]	add_u582;
wire		or_u1228_u0;
wire		and_u4105_u0;
reg		reg_20beb1e1_u0=1'h0;
wire	[15:0]	add_u583;
reg	[15:0]	syncEnable_u814_u0=16'h0;
wire		and_u4106_u0;
wire	[15:0]	mux_u426_u0;
wire	[15:0]	latch_02bc9e11_out;
reg	[15:0]	latch_02bc9e11_reg=16'h0;
wire		or_u1229_u0;
reg	[15:0]	syncEnable_u815_u0=16'h0;
reg		reg_1490018b_u0=1'h0;
assign simplePinWrite=GO&{1{GO}};
assign lessThanEqualTo_a_signed={mux_u425[15], mux_u425};
assign lessThanEqualTo_b_signed=17'h7;
assign lessThanEqualTo=lessThanEqualTo_a_signed<=lessThanEqualTo_b_signed;
assign and_u4097_u0=or_u1227_u0&not_u654_u0;
assign not_u654_u0=~lessThanEqualTo;
assign and_u4098_u0=or_u1227_u0&lessThanEqualTo;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_4a35a071_u0<=1'h0;
else reg_4a35a071_u0<=and_u4099_u0;
end
assign and_u4099_u0=and_u4098_u0&or_u1227_u0;
assign and_u4100_u0=and_u4097_u0&or_u1227_u0;
assign add={13'b0, port_7ee25a17_, 3'b0}+{mux_u425[15], mux_u425[15], mux_u425[15], mux_u425[15], mux_u425[15], mux_u425[15], mux_u425[15], mux_u425[15], mux_u425[15], mux_u425[15], mux_u425[15], mux_u425[15], mux_u425[15], mux_u425[15], mux_u425[15], mux_u425[15], mux_u425};
assign add_u579={add[20], add[20], add[20], add[20], add[20], add[20], add[20], add[20], add[20], add[20], add[20], add[20:0]}+32'h0;
always @(posedge CLK or posedge and_u4099_u0 or posedge or_u1226_u0)
begin
if (or_u1226_u0)
reg_6d0dbf08_u0<=1'h0;
else if (and_u4099_u0)
reg_6d0dbf08_u0<=1'h1;
else reg_6d0dbf08_u0<=reg_6d0dbf08_u0;
end
assign and_u4101_u0=reg_6d0dbf08_u0&port_4bf12c4e_;
assign or_u1226_u0=and_u4101_u0|RESET;
assign add_u580=mux_u425+16'h1;
always @(posedge CLK)
begin
if (and_u4099_u0)
syncEnable_u813<=add_u580;
end
assign mux_u425=(GO)?16'h0:syncEnable_u813;
assign or_u1227_u0=GO|reg_4a35a071_u0;
assign latch_43b8c804_out=(GO)?port_0266fa2c_:latch_43b8c804_reg;
always @(posedge CLK)
begin
if (GO)
latch_43b8c804_reg<=port_0266fa2c_;
end
assign add_u581=port_7ee25a17_+16'h1;
assign and_u4102_u0=and_u4103_u0&or_u1229_u0;
assign lessThanEqualTo_u5_a_signed={mux_u426_u0[15], mux_u426_u0};
assign lessThanEqualTo_u5_b_signed=17'h8;
assign lessThanEqualTo_u5=lessThanEqualTo_u5_a_signed<=lessThanEqualTo_u5_b_signed;
assign and_u4103_u0=or_u1229_u0&lessThanEqualTo_u5;
assign not_u655_u0=~lessThanEqualTo_u5;
assign and_u4104_u0=or_u1229_u0&not_u655_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u279<=1'h0;
else and_delayed_u279<=and_u4102_u0;
end
assign subtract=mux_u426_u0-16'h1;
assign add_u582={subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract[15], subtract}+32'h0;
assign or_u1228_u0=and_u4105_u0|RESET;
assign and_u4105_u0=reg_20beb1e1_u0&port_00eaa84f_;
always @(posedge CLK or posedge and_u4102_u0 or posedge or_u1228_u0)
begin
if (or_u1228_u0)
reg_20beb1e1_u0<=1'h0;
else if (and_u4102_u0)
reg_20beb1e1_u0<=1'h1;
else reg_20beb1e1_u0<=reg_20beb1e1_u0;
end
assign add_u583=mux_u426_u0+16'h1;
always @(posedge CLK)
begin
if (and_u4102_u0)
syncEnable_u814_u0<=add_u583;
end
assign and_u4106_u0=and_u4104_u0&or_u1229_u0;
assign mux_u426_u0=(GO)?16'h1:syncEnable_u814_u0;
assign latch_02bc9e11_out=(GO)?port_0266fa2c_:latch_02bc9e11_reg;
always @(posedge CLK)
begin
if (GO)
latch_02bc9e11_reg<=port_0266fa2c_;
end
assign or_u1229_u0=GO|and_delayed_u279;
always @(posedge CLK)
begin
if (GO)
syncEnable_u815_u0<=add_u581;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_1490018b_u0<=1'h0;
else reg_1490018b_u0<=and_u4100_u0;
end
assign RESULT=and_u4100_u0;
assign RESULT_u2399=syncEnable_u815_u0;
assign RESULT_u2400=and_u4102_u0;
assign RESULT_u2401=add_u582;
assign RESULT_u2402=latch_02bc9e11_out;
assign RESULT_u2403=3'h1;
assign RESULT_u2404=and_u4099_u0;
assign RESULT_u2405=add_u579;
assign RESULT_u2406=latch_43b8c804_out;
assign RESULT_u2407=3'h1;
assign RESULT_u2408=simplePinWrite;
assign DONE=reg_1490018b_u0;
endmodule



module resized_LH3_xy_structuralmemory_46badd45_(CLK_u24, bus_568ab95c_, bus_12817703_, bus_12f2a754_, bus_1cfe3bb9_, bus_183866fe_, bus_6170e247_, bus_04fa5f53_, bus_2186a09b_);
input		CLK_u24;
input		bus_568ab95c_;
input	[31:0]	bus_12817703_;
input	[2:0]	bus_12f2a754_;
input		bus_1cfe3bb9_;
input		bus_183866fe_;
input	[15:0]	bus_6170e247_;
output	[15:0]	bus_04fa5f53_;
output		bus_2186a09b_;
reg		logicalMem_47fabf37_we_delay0_u0=1'h0;
wire		and_6f46b1a7_u0;
wire		not_330a968c_u0;
wire		or_228946a0_u0;
wire		or_42d43119_u0;
wire	[15:0]	bus_3410ff1c_;
always @(posedge CLK_u24 or posedge bus_568ab95c_)
begin
if (bus_568ab95c_)
logicalMem_47fabf37_we_delay0_u0<=1'h0;
else logicalMem_47fabf37_we_delay0_u0<=bus_183866fe_;
end
assign and_6f46b1a7_u0=bus_1cfe3bb9_&not_330a968c_u0;
assign not_330a968c_u0=~bus_183866fe_;
assign or_228946a0_u0=and_6f46b1a7_u0|logicalMem_47fabf37_we_delay0_u0;
assign bus_04fa5f53_=bus_3410ff1c_;
assign bus_2186a09b_=or_228946a0_u0;
assign or_42d43119_u0=bus_1cfe3bb9_|bus_183866fe_;
resized_LH3_xy_forge_memory_512x16_43 resized_LH3_xy_forge_memory_512x16_43_instance1(.CLK(CLK_u24), 
  .EN(or_42d43119_u0), .WE(bus_183866fe_), .ADDR(bus_12817703_), .DIN(bus_6170e247_), 
  .DOUT(bus_3410ff1c_), .DONE());
endmodule


